// nios2.v

// Generated using ACDS version 13.0 156 at 2018.05.02.19:47:15

`timescale 1 ps / 1 ps
module nios2 (
		input  wire        clk_clk,                              //                  clk.clk
		input  wire        reset_reset_n,                        //                reset.reset_n
		output wire [0:0]  ddr2_mem_odt,                         //                 ddr2.mem_odt
		inout  wire [0:0]  ddr2_mem_clk,                         //                     .mem_clk
		inout  wire [0:0]  ddr2_mem_clk_n,                       //                     .mem_clk_n
		output wire [0:0]  ddr2_mem_cs_n,                        //                     .mem_cs_n
		output wire [0:0]  ddr2_mem_cke,                         //                     .mem_cke
		output wire [12:0] ddr2_mem_addr,                        //                     .mem_addr
		output wire [1:0]  ddr2_mem_ba,                          //                     .mem_ba
		output wire        ddr2_mem_ras_n,                       //                     .mem_ras_n
		output wire        ddr2_mem_cas_n,                       //                     .mem_cas_n
		output wire        ddr2_mem_we_n,                        //                     .mem_we_n
		inout  wire [15:0] ddr2_mem_dq,                          //                     .mem_dq
		inout  wire [1:0]  ddr2_mem_dqs,                         //                     .mem_dqs
		output wire [1:0]  ddr2_mem_dm,                          //                     .mem_dm
		output wire [5:0]  led_export,                           //                  led.export
		input  wire [3:0]  key_export,                           //                  key.export
		input  wire        uart_rxd,                             //                 uart.rxd
		output wire        uart_txd,                             //                     .txd
		input  wire        spi_dp_MISO,                          //               spi_dp.MISO
		output wire        spi_dp_MOSI,                          //                     .MOSI
		output wire        spi_dp_SCLK,                          //                     .SCLK
		output wire        spi_dp_SS_n,                          //                     .SS_n
		output wire        epcs_flash_dclk,                      //           epcs_flash.dclk
		output wire        epcs_flash_sce,                       //                     .sce
		output wire        epcs_flash_sdo,                       //                     .sdo
		input  wire        epcs_flash_data0,                     //                     .data0
		input  wire        spi_ad5781_MISO,                      //           spi_ad5781.MISO
		output wire        spi_ad5781_MOSI,                      //                     .MOSI
		output wire        spi_ad5781_SCLK,                      //                     .SCLK
		output wire        spi_ad5781_SS_n,                      //                     .SS_n
		output wire        nios_clk_clk,                         //             nios_clk.clk
		input  wire [13:0] ad9245_2_ad_data_export,              //     ad9245_2_ad_data.export
		input  wire [13:0] ad9245_1_ad_data_export,              //     ad9245_1_ad_data.export
		inout  wire        oc_i2c_master_scl_pad_io,             //        oc_i2c_master.scl_pad_io
		inout  wire        oc_i2c_master_sda_pad_io,             //                     .sda_pad_io
		input  wire        spi_master_miso,                      //           spi_master.miso
		output wire        spi_master_mosi,                      //                     .mosi
		output wire        spi_master_sclk,                      //                     .sclk
		output wire [0:0]  spi_master_ss,                        //                     .ss
		input  wire        ad9266_MISO,                          //               ad9266.MISO
		output wire        ad9266_MOSI,                          //                     .MOSI
		output wire        ad9266_SCLK,                          //                     .SCLK
		output wire        ad9266_SS_n,                          //                     .SS_n
		output wire [7:0]  clk_gen_clk_out_export,               //      clk_gen_clk_out.export
		output wire [13:0] dac2904_1_dac_data_export,            //   dac2904_1_dac_data.export
		input  wire        dac2904_1_sample_clk_clk,             // dac2904_1_sample_clk.clk
		output wire [13:0] dac2904_2_dac_data_export,            //   dac2904_2_dac_data.export
		input  wire        dac2904_2_sample_clk_clk,             // dac2904_2_sample_clk.clk
		output wire [13:0] dac2904_3_dac_data_export,            //   dac2904_3_dac_data.export
		input  wire        dac2904_3_sample_clk_clk,             // dac2904_3_sample_clk.clk
		output wire [13:0] dac2904_4_dac_data_export,            //   dac2904_4_dac_data.export
		input  wire        dac2904_4_sample_clk_clk,             // dac2904_4_sample_clk.clk
		output wire [13:0] wave_gen_0_dac_export,                //       wave_gen_0_dac.export
		output wire [13:0] demodulation_0_ad_da_dac,             // demodulation_0_ad_da.dac
		input  wire [13:0] demodulation_0_ad_da_ad,              //                     .ad
		input  wire        demodulation_0_ad_da_modulation_wave, //                     .modulation_wave
		output wire [13:0] wave_gen_1_dac_export,                //       wave_gen_1_dac.export
		output wire [13:0] wave_gen_2_dac_export                 //       wave_gen_2_dac.export
	);

	wire          altpll_0_c0_clk;                                                                                    // altpll_0:c0 -> [ad9245_1:clk, ad9245_1_s1_translator:clk, ad9245_1_s1_translator_avalon_universal_slave_0_agent:clk, ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, ad9245_2:clk, ad9245_2_s1_translator:clk, ad9245_2_s1_translator_avalon_universal_slave_0_agent:clk, ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, ad9266:clk, ad9266_spi_control_port_translator:clk, ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:clk, ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router_003:clk, clk_gen:clk, clk_gen_s1_translator:clk, clk_gen_s1_translator_avalon_universal_slave_0_agent:clk, clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux_003:clk, cmd_xbar_mux_021:clk, cmd_xbar_mux_022:clk, crosser:in_clk, crosser_001:out_clk, crosser_002:out_clk, crosser_003:out_clk, crosser_004:in_clk, crosser_005:in_clk, dac2904_1:clk, dac2904_1_s0_translator:clk, dac2904_1_s0_translator_avalon_universal_slave_0_agent:clk, dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, dac2904_2:clk, dac2904_2_s0_translator:clk, dac2904_2_s0_translator_avalon_universal_slave_0_agent:clk, dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, dac2904_3:clk, dac2904_3_s0_translator:clk, dac2904_3_s0_translator_avalon_universal_slave_0_agent:clk, dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, dac2904_4:clk, dac2904_4_s0_translator:clk, dac2904_4_s0_translator_avalon_universal_slave_0_agent:clk, dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, demodulation_0:clk, demodulation_0_s0_translator:clk, demodulation_0_s0_translator_avalon_universal_slave_0_agent:clk, demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, id_router_016:clk, id_router_017:clk, id_router_018:clk, id_router_019:clk, id_router_020:clk, id_router_021:clk, id_router_022:clk, id_router_023:clk, id_router_024:clk, id_router_025:clk, id_router_026:clk, id_router_027:clk, id_router_028:clk, id_router_029:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_002:receiver_clk, irq_synchronizer_003:receiver_clk, irq_synchronizer_004:receiver_clk, irq_synchronizer_005:receiver_clk, irq_synchronizer_006:receiver_clk, irq_synchronizer_007:receiver_clk, irq_synchronizer_008:receiver_clk, irq_synchronizer_009:receiver_clk, jtag_uart_0:clk, jtag_uart_0_avalon_jtag_slave_translator:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter_001:clk, oc_i2c_master_0:wb_clk_i, oc_i2c_master_0_s1_translator:clk, oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:clk, oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_key:clk, pio_key_s1_translator:clk, pio_key_s1_translator_avalon_universal_slave_0_agent:clk, pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_led:clk, pio_led_s1_translator:clk, pio_led_s1_translator_avalon_universal_slave_0_agent:clk, pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_demux_016:clk, rsp_xbar_demux_017:clk, rsp_xbar_demux_018:clk, rsp_xbar_demux_019:clk, rsp_xbar_demux_020:clk, rsp_xbar_demux_021:clk, rsp_xbar_demux_022:clk, rsp_xbar_demux_023:clk, rsp_xbar_demux_024:clk, rsp_xbar_demux_025:clk, rsp_xbar_demux_026:clk, rsp_xbar_demux_027:clk, rsp_xbar_demux_028:clk, rsp_xbar_demux_029:clk, rsp_xbar_mux_003:clk, rst_controller_001:clk, slow_peripheral_bridge:m0_clk, slow_peripheral_bridge_m0_translator:clk, slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:clk, spi_0:clk, spi_0_spi_control_port_translator:clk, spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:clk, spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, spi_ad5781:clk, spi_ad5781_spi_control_port_translator:clk, spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:clk, spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, spi_master_0:clk, spi_master_0_s1_translator:clk, spi_master_0_s1_translator_avalon_universal_slave_0_agent:clk, spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sysid:clock, sysid_control_slave_translator:clk, sysid_control_slave_translator_avalon_universal_slave_0_agent:clk, sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, systimer:clk, systimer_s1_translator:clk, systimer_s1_translator_avalon_universal_slave_0_agent:clk, systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timestamp:clk, timestamp_s1_translator:clk, timestamp_s1_translator_avalon_universal_slave_0_agent:clk, timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, uart_0:clk, uart_0_s1_translator:clk, uart_0_s1_translator_avalon_universal_slave_0_agent:clk, uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, wave_gen_0:clk, wave_gen_0_s0_translator:clk, wave_gen_0_s0_translator_avalon_universal_slave_0_agent:clk, wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, wave_gen_1:clk, wave_gen_1_s0_translator:clk, wave_gen_1_s0_translator_avalon_universal_slave_0_agent:clk, wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, wave_gen_2:clk, wave_gen_2_s0_translator:clk, wave_gen_2_s0_translator_avalon_universal_slave_0_agent:clk, wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk]
	wire          ddr2_sysclk_clk;                                                                                    // ddr2:phy_clk -> [addr_router_005:clk, cmd_xbar_demux_005:clk, cpu_ddr2_clock_bridge:m0_clk, cpu_ddr2_clock_bridge_m0_translator:clk, cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:clk, ddr2_s1_translator:clk, ddr2_s1_translator_avalon_universal_slave_0_agent:clk, ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router_030:clk, rsp_xbar_demux_030:clk, rst_controller_005:clk]
	wire          altpll_0_c1_clk;                                                                                    // altpll_0:c1 -> [ddr2:pll_ref_clk, rst_controller_002:clk, rst_controller_003:clk]
	wire          nios2_instruction_master_waitrequest;                                                               // nios2_instruction_master_translator:av_waitrequest -> nios2:i_waitrequest
	wire   [26:0] nios2_instruction_master_address;                                                                   // nios2:i_address -> nios2_instruction_master_translator:av_address
	wire          nios2_instruction_master_read;                                                                      // nios2:i_read -> nios2_instruction_master_translator:av_read
	wire   [31:0] nios2_instruction_master_readdata;                                                                  // nios2_instruction_master_translator:av_readdata -> nios2:i_readdata
	wire          nios2_instruction_master_readdatavalid;                                                             // nios2_instruction_master_translator:av_readdatavalid -> nios2:i_readdatavalid
	wire          nios2_data_master_waitrequest;                                                                      // nios2_data_master_translator:av_waitrequest -> nios2:d_waitrequest
	wire   [31:0] nios2_data_master_writedata;                                                                        // nios2:d_writedata -> nios2_data_master_translator:av_writedata
	wire   [26:0] nios2_data_master_address;                                                                          // nios2:d_address -> nios2_data_master_translator:av_address
	wire          nios2_data_master_write;                                                                            // nios2:d_write -> nios2_data_master_translator:av_write
	wire          nios2_data_master_read;                                                                             // nios2:d_read -> nios2_data_master_translator:av_read
	wire   [31:0] nios2_data_master_readdata;                                                                         // nios2_data_master_translator:av_readdata -> nios2:d_readdata
	wire          nios2_data_master_debugaccess;                                                                      // nios2:jtag_debug_module_debugaccess_to_roms -> nios2_data_master_translator:av_debugaccess
	wire    [3:0] nios2_data_master_byteenable;                                                                       // nios2:d_byteenable -> nios2_data_master_translator:av_byteenable
	wire          dma_0_read_master_waitrequest;                                                                      // dma_0_read_master_translator:av_waitrequest -> dma_0:read_waitrequest
	wire   [26:0] dma_0_read_master_address;                                                                          // dma_0:read_address -> dma_0_read_master_translator:av_address
	wire          dma_0_read_master_chipselect;                                                                       // dma_0:read_chipselect -> dma_0_read_master_translator:av_chipselect
	wire          dma_0_read_master_read;                                                                             // dma_0:read_read_n -> dma_0_read_master_translator:av_read
	wire   [31:0] dma_0_read_master_readdata;                                                                         // dma_0_read_master_translator:av_readdata -> dma_0:read_readdata
	wire          dma_0_read_master_readdatavalid;                                                                    // dma_0_read_master_translator:av_readdatavalid -> dma_0:read_readdatavalid
	wire          nios2_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                 // nios2:jtag_debug_module_waitrequest -> nios2_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // nios2_jtag_debug_module_translator:av_writedata -> nios2:jtag_debug_module_writedata
	wire    [8:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // nios2_jtag_debug_module_translator:av_address -> nios2:jtag_debug_module_address
	wire          nios2_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // nios2_jtag_debug_module_translator:av_write -> nios2:jtag_debug_module_write
	wire          nios2_jtag_debug_module_translator_avalon_anti_slave_0_read;                                        // nios2_jtag_debug_module_translator:av_read -> nios2:jtag_debug_module_read
	wire   [31:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // nios2:jtag_debug_module_readdata -> nios2_jtag_debug_module_translator:av_readdata
	wire          nios2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // nios2_jtag_debug_module_translator:av_debugaccess -> nios2:jtag_debug_module_debugaccess
	wire    [3:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // nios2_jtag_debug_module_translator:av_byteenable -> nios2:jtag_debug_module_byteenable
	wire   [31:0] epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_writedata;                              // epcs_flash_epcs_control_port_translator:av_writedata -> epcs_flash:writedata
	wire    [8:0] epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_address;                                // epcs_flash_epcs_control_port_translator:av_address -> epcs_flash:address
	wire          epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_chipselect;                             // epcs_flash_epcs_control_port_translator:av_chipselect -> epcs_flash:chipselect
	wire          epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_write;                                  // epcs_flash_epcs_control_port_translator:av_write -> epcs_flash:write_n
	wire          epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_read;                                   // epcs_flash_epcs_control_port_translator:av_read -> epcs_flash:read_n
	wire   [31:0] epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_readdata;                               // epcs_flash:readdata -> epcs_flash_epcs_control_port_translator:av_readdata
	wire   [31:0] onchip_ram_s1_translator_avalon_anti_slave_0_writedata;                                             // onchip_ram_s1_translator:av_writedata -> onchip_ram:writedata
	wire    [9:0] onchip_ram_s1_translator_avalon_anti_slave_0_address;                                               // onchip_ram_s1_translator:av_address -> onchip_ram:address
	wire          onchip_ram_s1_translator_avalon_anti_slave_0_chipselect;                                            // onchip_ram_s1_translator:av_chipselect -> onchip_ram:chipselect
	wire          onchip_ram_s1_translator_avalon_anti_slave_0_clken;                                                 // onchip_ram_s1_translator:av_clken -> onchip_ram:clken
	wire          onchip_ram_s1_translator_avalon_anti_slave_0_write;                                                 // onchip_ram_s1_translator:av_write -> onchip_ram:write
	wire   [31:0] onchip_ram_s1_translator_avalon_anti_slave_0_readdata;                                              // onchip_ram:readdata -> onchip_ram_s1_translator:av_readdata
	wire    [3:0] onchip_ram_s1_translator_avalon_anti_slave_0_byteenable;                                            // onchip_ram_s1_translator:av_byteenable -> onchip_ram:byteenable
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                // cpu_ddr2_clock_bridge:s0_waitrequest -> cpu_ddr2_clock_bridge_s0_translator:av_waitrequest
	wire    [0:0] cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount;                                 // cpu_ddr2_clock_bridge_s0_translator:av_burstcount -> cpu_ddr2_clock_bridge:s0_burstcount
	wire   [31:0] cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_writedata;                                  // cpu_ddr2_clock_bridge_s0_translator:av_writedata -> cpu_ddr2_clock_bridge:s0_writedata
	wire   [25:0] cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_address;                                    // cpu_ddr2_clock_bridge_s0_translator:av_address -> cpu_ddr2_clock_bridge:s0_address
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_write;                                      // cpu_ddr2_clock_bridge_s0_translator:av_write -> cpu_ddr2_clock_bridge:s0_write
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_read;                                       // cpu_ddr2_clock_bridge_s0_translator:av_read -> cpu_ddr2_clock_bridge:s0_read
	wire   [31:0] cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_readdata;                                   // cpu_ddr2_clock_bridge:s0_readdata -> cpu_ddr2_clock_bridge_s0_translator:av_readdata
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                                // cpu_ddr2_clock_bridge_s0_translator:av_debugaccess -> cpu_ddr2_clock_bridge:s0_debugaccess
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                              // cpu_ddr2_clock_bridge:s0_readdatavalid -> cpu_ddr2_clock_bridge_s0_translator:av_readdatavalid
	wire    [3:0] cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable;                                 // cpu_ddr2_clock_bridge_s0_translator:av_byteenable -> cpu_ddr2_clock_bridge:s0_byteenable
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                               // slow_peripheral_bridge:s0_waitrequest -> slow_peripheral_bridge_s0_translator:av_waitrequest
	wire    [0:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount;                                // slow_peripheral_bridge_s0_translator:av_burstcount -> slow_peripheral_bridge:s0_burstcount
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata;                                 // slow_peripheral_bridge_s0_translator:av_writedata -> slow_peripheral_bridge:s0_writedata
	wire    [9:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_address;                                   // slow_peripheral_bridge_s0_translator:av_address -> slow_peripheral_bridge:s0_address
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_write;                                     // slow_peripheral_bridge_s0_translator:av_write -> slow_peripheral_bridge:s0_write
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_read;                                      // slow_peripheral_bridge_s0_translator:av_read -> slow_peripheral_bridge:s0_read
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata;                                  // slow_peripheral_bridge:s0_readdata -> slow_peripheral_bridge_s0_translator:av_readdata
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                               // slow_peripheral_bridge_s0_translator:av_debugaccess -> slow_peripheral_bridge:s0_debugaccess
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                             // slow_peripheral_bridge:s0_readdatavalid -> slow_peripheral_bridge_s0_translator:av_readdatavalid
	wire    [3:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable;                                // slow_peripheral_bridge_s0_translator:av_byteenable -> slow_peripheral_bridge:s0_byteenable
	wire   [26:0] dma_0_control_port_slave_translator_avalon_anti_slave_0_writedata;                                  // dma_0_control_port_slave_translator:av_writedata -> dma_0:dma_ctl_writedata
	wire    [2:0] dma_0_control_port_slave_translator_avalon_anti_slave_0_address;                                    // dma_0_control_port_slave_translator:av_address -> dma_0:dma_ctl_address
	wire          dma_0_control_port_slave_translator_avalon_anti_slave_0_chipselect;                                 // dma_0_control_port_slave_translator:av_chipselect -> dma_0:dma_ctl_chipselect
	wire          dma_0_control_port_slave_translator_avalon_anti_slave_0_write;                                      // dma_0_control_port_slave_translator:av_write -> dma_0:dma_ctl_write_n
	wire   [26:0] dma_0_control_port_slave_translator_avalon_anti_slave_0_readdata;                                   // dma_0:dma_ctl_readdata -> dma_0_control_port_slave_translator:av_readdata
	wire    [0:0] slow_peripheral_bridge_m0_burstcount;                                                               // slow_peripheral_bridge:m0_burstcount -> slow_peripheral_bridge_m0_translator:av_burstcount
	wire          slow_peripheral_bridge_m0_waitrequest;                                                              // slow_peripheral_bridge_m0_translator:av_waitrequest -> slow_peripheral_bridge:m0_waitrequest
	wire    [9:0] slow_peripheral_bridge_m0_address;                                                                  // slow_peripheral_bridge:m0_address -> slow_peripheral_bridge_m0_translator:av_address
	wire   [31:0] slow_peripheral_bridge_m0_writedata;                                                                // slow_peripheral_bridge:m0_writedata -> slow_peripheral_bridge_m0_translator:av_writedata
	wire          slow_peripheral_bridge_m0_write;                                                                    // slow_peripheral_bridge:m0_write -> slow_peripheral_bridge_m0_translator:av_write
	wire          slow_peripheral_bridge_m0_read;                                                                     // slow_peripheral_bridge:m0_read -> slow_peripheral_bridge_m0_translator:av_read
	wire   [31:0] slow_peripheral_bridge_m0_readdata;                                                                 // slow_peripheral_bridge_m0_translator:av_readdata -> slow_peripheral_bridge:m0_readdata
	wire          slow_peripheral_bridge_m0_debugaccess;                                                              // slow_peripheral_bridge:m0_debugaccess -> slow_peripheral_bridge_m0_translator:av_debugaccess
	wire    [3:0] slow_peripheral_bridge_m0_byteenable;                                                               // slow_peripheral_bridge:m0_byteenable -> slow_peripheral_bridge_m0_translator:av_byteenable
	wire          slow_peripheral_bridge_m0_readdatavalid;                                                            // slow_peripheral_bridge_m0_translator:av_readdatavalid -> slow_peripheral_bridge:m0_readdatavalid
	wire          dma_0_write_master_waitrequest;                                                                     // dma_0_write_master_translator:av_waitrequest -> dma_0:write_waitrequest
	wire   [31:0] dma_0_write_master_writedata;                                                                       // dma_0:write_writedata -> dma_0_write_master_translator:av_writedata
	wire    [9:0] dma_0_write_master_address;                                                                         // dma_0:write_address -> dma_0_write_master_translator:av_address
	wire          dma_0_write_master_chipselect;                                                                      // dma_0:write_chipselect -> dma_0_write_master_translator:av_chipselect
	wire          dma_0_write_master_write;                                                                           // dma_0:write_write_n -> dma_0_write_master_translator:av_write
	wire    [3:0] dma_0_write_master_byteenable;                                                                      // dma_0:write_byteenable -> dma_0_write_master_translator:av_byteenable
	wire   [31:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata;                                        // altpll_0_pll_slave_translator:av_writedata -> altpll_0:writedata
	wire    [1:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_address;                                          // altpll_0_pll_slave_translator:av_address -> altpll_0:address
	wire          altpll_0_pll_slave_translator_avalon_anti_slave_0_write;                                            // altpll_0_pll_slave_translator:av_write -> altpll_0:write
	wire          altpll_0_pll_slave_translator_avalon_anti_slave_0_read;                                             // altpll_0_pll_slave_translator:av_read -> altpll_0:read
	wire   [31:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata;                                         // altpll_0:readdata -> altpll_0_pll_slave_translator:av_readdata
	wire    [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                         // sysid_control_slave_translator:av_address -> sysid:address
	wire   [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                        // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire    [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] systimer_s1_translator_avalon_anti_slave_0_writedata;                                               // systimer_s1_translator:av_writedata -> systimer:writedata
	wire    [2:0] systimer_s1_translator_avalon_anti_slave_0_address;                                                 // systimer_s1_translator:av_address -> systimer:address
	wire          systimer_s1_translator_avalon_anti_slave_0_chipselect;                                              // systimer_s1_translator:av_chipselect -> systimer:chipselect
	wire          systimer_s1_translator_avalon_anti_slave_0_write;                                                   // systimer_s1_translator:av_write -> systimer:write_n
	wire   [15:0] systimer_s1_translator_avalon_anti_slave_0_readdata;                                                // systimer:readdata -> systimer_s1_translator:av_readdata
	wire   [31:0] pio_key_s1_translator_avalon_anti_slave_0_writedata;                                                // pio_key_s1_translator:av_writedata -> pio_key:writedata
	wire    [1:0] pio_key_s1_translator_avalon_anti_slave_0_address;                                                  // pio_key_s1_translator:av_address -> pio_key:address
	wire          pio_key_s1_translator_avalon_anti_slave_0_chipselect;                                               // pio_key_s1_translator:av_chipselect -> pio_key:chipselect
	wire          pio_key_s1_translator_avalon_anti_slave_0_write;                                                    // pio_key_s1_translator:av_write -> pio_key:write_n
	wire   [31:0] pio_key_s1_translator_avalon_anti_slave_0_readdata;                                                 // pio_key:readdata -> pio_key_s1_translator:av_readdata
	wire   [15:0] spi_0_spi_control_port_translator_avalon_anti_slave_0_writedata;                                    // spi_0_spi_control_port_translator:av_writedata -> spi_0:data_from_cpu
	wire    [2:0] spi_0_spi_control_port_translator_avalon_anti_slave_0_address;                                      // spi_0_spi_control_port_translator:av_address -> spi_0:mem_addr
	wire          spi_0_spi_control_port_translator_avalon_anti_slave_0_chipselect;                                   // spi_0_spi_control_port_translator:av_chipselect -> spi_0:spi_select
	wire          spi_0_spi_control_port_translator_avalon_anti_slave_0_write;                                        // spi_0_spi_control_port_translator:av_write -> spi_0:write_n
	wire          spi_0_spi_control_port_translator_avalon_anti_slave_0_read;                                         // spi_0_spi_control_port_translator:av_read -> spi_0:read_n
	wire   [15:0] spi_0_spi_control_port_translator_avalon_anti_slave_0_readdata;                                     // spi_0:data_to_cpu -> spi_0_spi_control_port_translator:av_readdata
	wire   [15:0] uart_0_s1_translator_avalon_anti_slave_0_writedata;                                                 // uart_0_s1_translator:av_writedata -> uart_0:writedata
	wire    [2:0] uart_0_s1_translator_avalon_anti_slave_0_address;                                                   // uart_0_s1_translator:av_address -> uart_0:address
	wire          uart_0_s1_translator_avalon_anti_slave_0_chipselect;                                                // uart_0_s1_translator:av_chipselect -> uart_0:chipselect
	wire          uart_0_s1_translator_avalon_anti_slave_0_write;                                                     // uart_0_s1_translator:av_write -> uart_0:write_n
	wire          uart_0_s1_translator_avalon_anti_slave_0_read;                                                      // uart_0_s1_translator:av_read -> uart_0:read_n
	wire   [15:0] uart_0_s1_translator_avalon_anti_slave_0_readdata;                                                  // uart_0:readdata -> uart_0_s1_translator:av_readdata
	wire          uart_0_s1_translator_avalon_anti_slave_0_begintransfer;                                             // uart_0_s1_translator:av_begintransfer -> uart_0:begintransfer
	wire   [31:0] pio_led_s1_translator_avalon_anti_slave_0_writedata;                                                // pio_led_s1_translator:av_writedata -> pio_led:writedata
	wire    [1:0] pio_led_s1_translator_avalon_anti_slave_0_address;                                                  // pio_led_s1_translator:av_address -> pio_led:address
	wire          pio_led_s1_translator_avalon_anti_slave_0_chipselect;                                               // pio_led_s1_translator:av_chipselect -> pio_led:chipselect
	wire          pio_led_s1_translator_avalon_anti_slave_0_write;                                                    // pio_led_s1_translator:av_write -> pio_led:write_n
	wire   [31:0] pio_led_s1_translator_avalon_anti_slave_0_readdata;                                                 // pio_led:readdata -> pio_led_s1_translator:av_readdata
	wire   [15:0] timestamp_s1_translator_avalon_anti_slave_0_writedata;                                              // timestamp_s1_translator:av_writedata -> timestamp:writedata
	wire    [2:0] timestamp_s1_translator_avalon_anti_slave_0_address;                                                // timestamp_s1_translator:av_address -> timestamp:address
	wire          timestamp_s1_translator_avalon_anti_slave_0_chipselect;                                             // timestamp_s1_translator:av_chipselect -> timestamp:chipselect
	wire          timestamp_s1_translator_avalon_anti_slave_0_write;                                                  // timestamp_s1_translator:av_write -> timestamp:write_n
	wire   [15:0] timestamp_s1_translator_avalon_anti_slave_0_readdata;                                               // timestamp:readdata -> timestamp_s1_translator:av_readdata
	wire   [15:0] spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_writedata;                               // spi_ad5781_spi_control_port_translator:av_writedata -> spi_ad5781:data_from_cpu
	wire    [2:0] spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_address;                                 // spi_ad5781_spi_control_port_translator:av_address -> spi_ad5781:mem_addr
	wire          spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_chipselect;                              // spi_ad5781_spi_control_port_translator:av_chipselect -> spi_ad5781:spi_select
	wire          spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_write;                                   // spi_ad5781_spi_control_port_translator:av_write -> spi_ad5781:write_n
	wire          spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_read;                                    // spi_ad5781_spi_control_port_translator:av_read -> spi_ad5781:read_n
	wire   [15:0] spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_readdata;                                // spi_ad5781:data_to_cpu -> spi_ad5781_spi_control_port_translator:av_readdata
	wire          ad9245_2_s1_translator_avalon_anti_slave_0_chipselect;                                              // ad9245_2_s1_translator:av_chipselect -> ad9245_2:chipselect
	wire          ad9245_2_s1_translator_avalon_anti_slave_0_read;                                                    // ad9245_2_s1_translator:av_read -> ad9245_2:read
	wire   [31:0] ad9245_2_s1_translator_avalon_anti_slave_0_readdata;                                                // ad9245_2:readdata -> ad9245_2_s1_translator:av_readdata
	wire   [31:0] clk_gen_s1_translator_avalon_anti_slave_0_writedata;                                                // clk_gen_s1_translator:av_writedata -> clk_gen:writedata
	wire    [4:0] clk_gen_s1_translator_avalon_anti_slave_0_address;                                                  // clk_gen_s1_translator:av_address -> clk_gen:address
	wire          clk_gen_s1_translator_avalon_anti_slave_0_chipselect;                                               // clk_gen_s1_translator:av_chipselect -> clk_gen:chipselect
	wire          clk_gen_s1_translator_avalon_anti_slave_0_write;                                                    // clk_gen_s1_translator:av_write -> clk_gen:write
	wire          clk_gen_s1_translator_avalon_anti_slave_0_read;                                                     // clk_gen_s1_translator:av_read -> clk_gen:read
	wire   [31:0] clk_gen_s1_translator_avalon_anti_slave_0_readdata;                                                 // clk_gen:readdata -> clk_gen_s1_translator:av_readdata
	wire          oc_i2c_master_0_s1_translator_avalon_anti_slave_0_waitrequest;                                      // oc_i2c_master_0:wb_ack_o -> oc_i2c_master_0_s1_translator:av_waitrequest
	wire   [31:0] oc_i2c_master_0_s1_translator_avalon_anti_slave_0_writedata;                                        // oc_i2c_master_0_s1_translator:av_writedata -> oc_i2c_master_0:wb_dat_i
	wire    [2:0] oc_i2c_master_0_s1_translator_avalon_anti_slave_0_address;                                          // oc_i2c_master_0_s1_translator:av_address -> oc_i2c_master_0:wb_adr_i
	wire          oc_i2c_master_0_s1_translator_avalon_anti_slave_0_chipselect;                                       // oc_i2c_master_0_s1_translator:av_chipselect -> oc_i2c_master_0:wb_cyc_i
	wire          oc_i2c_master_0_s1_translator_avalon_anti_slave_0_write;                                            // oc_i2c_master_0_s1_translator:av_write -> oc_i2c_master_0:wb_we_i
	wire   [31:0] oc_i2c_master_0_s1_translator_avalon_anti_slave_0_readdata;                                         // oc_i2c_master_0:wb_dat_o -> oc_i2c_master_0_s1_translator:av_readdata
	wire          oc_i2c_master_0_s1_translator_avalon_anti_slave_0_begintransfer;                                    // oc_i2c_master_0_s1_translator:av_begintransfer -> oc_i2c_master_0:wb_stb_i
	wire   [31:0] spi_master_0_s1_translator_avalon_anti_slave_0_writedata;                                           // spi_master_0_s1_translator:av_writedata -> spi_master_0:writedata
	wire    [2:0] spi_master_0_s1_translator_avalon_anti_slave_0_address;                                             // spi_master_0_s1_translator:av_address -> spi_master_0:address
	wire          spi_master_0_s1_translator_avalon_anti_slave_0_chipselect;                                          // spi_master_0_s1_translator:av_chipselect -> spi_master_0:chipselect
	wire          spi_master_0_s1_translator_avalon_anti_slave_0_write;                                               // spi_master_0_s1_translator:av_write -> spi_master_0:write
	wire          spi_master_0_s1_translator_avalon_anti_slave_0_read;                                                // spi_master_0_s1_translator:av_read -> spi_master_0:read
	wire   [31:0] spi_master_0_s1_translator_avalon_anti_slave_0_readdata;                                            // spi_master_0:readdata -> spi_master_0_s1_translator:av_readdata
	wire   [15:0] ad9266_spi_control_port_translator_avalon_anti_slave_0_writedata;                                   // ad9266_spi_control_port_translator:av_writedata -> ad9266:data_from_cpu
	wire    [2:0] ad9266_spi_control_port_translator_avalon_anti_slave_0_address;                                     // ad9266_spi_control_port_translator:av_address -> ad9266:mem_addr
	wire          ad9266_spi_control_port_translator_avalon_anti_slave_0_chipselect;                                  // ad9266_spi_control_port_translator:av_chipselect -> ad9266:spi_select
	wire          ad9266_spi_control_port_translator_avalon_anti_slave_0_write;                                       // ad9266_spi_control_port_translator:av_write -> ad9266:write_n
	wire          ad9266_spi_control_port_translator_avalon_anti_slave_0_read;                                        // ad9266_spi_control_port_translator:av_read -> ad9266:read_n
	wire   [15:0] ad9266_spi_control_port_translator_avalon_anti_slave_0_readdata;                                    // ad9266:data_to_cpu -> ad9266_spi_control_port_translator:av_readdata
	wire          ad9245_1_s1_translator_avalon_anti_slave_0_chipselect;                                              // ad9245_1_s1_translator:av_chipselect -> ad9245_1:chipselect
	wire          ad9245_1_s1_translator_avalon_anti_slave_0_read;                                                    // ad9245_1_s1_translator:av_read -> ad9245_1:read
	wire   [31:0] ad9245_1_s1_translator_avalon_anti_slave_0_readdata;                                                // ad9245_1:readdata -> ad9245_1_s1_translator:av_readdata
	wire          dac2904_1_s0_translator_avalon_anti_slave_0_waitrequest;                                            // dac2904_1:avs_s0_waitrequest -> dac2904_1_s0_translator:av_waitrequest
	wire   [31:0] dac2904_1_s0_translator_avalon_anti_slave_0_writedata;                                              // dac2904_1_s0_translator:av_writedata -> dac2904_1:avs_s0_writedata
	wire          dac2904_1_s0_translator_avalon_anti_slave_0_chipselect;                                             // dac2904_1_s0_translator:av_chipselect -> dac2904_1:avs_s0_chipselect
	wire          dac2904_1_s0_translator_avalon_anti_slave_0_write;                                                  // dac2904_1_s0_translator:av_write -> dac2904_1:avs_s0_write
	wire          dac2904_2_s0_translator_avalon_anti_slave_0_waitrequest;                                            // dac2904_2:avs_s0_waitrequest -> dac2904_2_s0_translator:av_waitrequest
	wire   [31:0] dac2904_2_s0_translator_avalon_anti_slave_0_writedata;                                              // dac2904_2_s0_translator:av_writedata -> dac2904_2:avs_s0_writedata
	wire          dac2904_2_s0_translator_avalon_anti_slave_0_chipselect;                                             // dac2904_2_s0_translator:av_chipselect -> dac2904_2:avs_s0_chipselect
	wire          dac2904_2_s0_translator_avalon_anti_slave_0_write;                                                  // dac2904_2_s0_translator:av_write -> dac2904_2:avs_s0_write
	wire          dac2904_3_s0_translator_avalon_anti_slave_0_waitrequest;                                            // dac2904_3:avs_s0_waitrequest -> dac2904_3_s0_translator:av_waitrequest
	wire   [31:0] dac2904_3_s0_translator_avalon_anti_slave_0_writedata;                                              // dac2904_3_s0_translator:av_writedata -> dac2904_3:avs_s0_writedata
	wire          dac2904_3_s0_translator_avalon_anti_slave_0_chipselect;                                             // dac2904_3_s0_translator:av_chipselect -> dac2904_3:avs_s0_chipselect
	wire          dac2904_3_s0_translator_avalon_anti_slave_0_write;                                                  // dac2904_3_s0_translator:av_write -> dac2904_3:avs_s0_write
	wire          dac2904_4_s0_translator_avalon_anti_slave_0_waitrequest;                                            // dac2904_4:avs_s0_waitrequest -> dac2904_4_s0_translator:av_waitrequest
	wire   [31:0] dac2904_4_s0_translator_avalon_anti_slave_0_writedata;                                              // dac2904_4_s0_translator:av_writedata -> dac2904_4:avs_s0_writedata
	wire          dac2904_4_s0_translator_avalon_anti_slave_0_chipselect;                                             // dac2904_4_s0_translator:av_chipselect -> dac2904_4:avs_s0_chipselect
	wire          dac2904_4_s0_translator_avalon_anti_slave_0_write;                                                  // dac2904_4_s0_translator:av_write -> dac2904_4:avs_s0_write
	wire   [31:0] wave_gen_0_s0_translator_avalon_anti_slave_0_writedata;                                             // wave_gen_0_s0_translator:av_writedata -> wave_gen_0:avs_s0_writedata
	wire    [2:0] wave_gen_0_s0_translator_avalon_anti_slave_0_address;                                               // wave_gen_0_s0_translator:av_address -> wave_gen_0:avs_s0_address
	wire          wave_gen_0_s0_translator_avalon_anti_slave_0_chipselect;                                            // wave_gen_0_s0_translator:av_chipselect -> wave_gen_0:avs_s0_chipselect
	wire          wave_gen_0_s0_translator_avalon_anti_slave_0_write;                                                 // wave_gen_0_s0_translator:av_write -> wave_gen_0:avs_s0_write
	wire          wave_gen_0_s0_translator_avalon_anti_slave_0_read;                                                  // wave_gen_0_s0_translator:av_read -> wave_gen_0:avs_s0_read
	wire   [31:0] wave_gen_0_s0_translator_avalon_anti_slave_0_readdata;                                              // wave_gen_0:avs_s0_readdata -> wave_gen_0_s0_translator:av_readdata
	wire   [31:0] demodulation_0_s0_translator_avalon_anti_slave_0_writedata;                                         // demodulation_0_s0_translator:av_writedata -> demodulation_0:avs_s0_writedata
	wire    [2:0] demodulation_0_s0_translator_avalon_anti_slave_0_address;                                           // demodulation_0_s0_translator:av_address -> demodulation_0:avs_s0_address
	wire          demodulation_0_s0_translator_avalon_anti_slave_0_chipselect;                                        // demodulation_0_s0_translator:av_chipselect -> demodulation_0:avs_s0_chipselect
	wire          demodulation_0_s0_translator_avalon_anti_slave_0_write;                                             // demodulation_0_s0_translator:av_write -> demodulation_0:avs_s0_write
	wire          demodulation_0_s0_translator_avalon_anti_slave_0_read;                                              // demodulation_0_s0_translator:av_read -> demodulation_0:avs_s0_read
	wire   [31:0] demodulation_0_s0_translator_avalon_anti_slave_0_readdata;                                          // demodulation_0:avs_s0_readdata -> demodulation_0_s0_translator:av_readdata
	wire   [31:0] wave_gen_1_s0_translator_avalon_anti_slave_0_writedata;                                             // wave_gen_1_s0_translator:av_writedata -> wave_gen_1:avs_s0_writedata
	wire    [2:0] wave_gen_1_s0_translator_avalon_anti_slave_0_address;                                               // wave_gen_1_s0_translator:av_address -> wave_gen_1:avs_s0_address
	wire          wave_gen_1_s0_translator_avalon_anti_slave_0_chipselect;                                            // wave_gen_1_s0_translator:av_chipselect -> wave_gen_1:avs_s0_chipselect
	wire          wave_gen_1_s0_translator_avalon_anti_slave_0_write;                                                 // wave_gen_1_s0_translator:av_write -> wave_gen_1:avs_s0_write
	wire          wave_gen_1_s0_translator_avalon_anti_slave_0_read;                                                  // wave_gen_1_s0_translator:av_read -> wave_gen_1:avs_s0_read
	wire   [31:0] wave_gen_1_s0_translator_avalon_anti_slave_0_readdata;                                              // wave_gen_1:avs_s0_readdata -> wave_gen_1_s0_translator:av_readdata
	wire   [31:0] wave_gen_2_s0_translator_avalon_anti_slave_0_writedata;                                             // wave_gen_2_s0_translator:av_writedata -> wave_gen_2:avs_s0_writedata
	wire    [2:0] wave_gen_2_s0_translator_avalon_anti_slave_0_address;                                               // wave_gen_2_s0_translator:av_address -> wave_gen_2:avs_s0_address
	wire          wave_gen_2_s0_translator_avalon_anti_slave_0_chipselect;                                            // wave_gen_2_s0_translator:av_chipselect -> wave_gen_2:avs_s0_chipselect
	wire          wave_gen_2_s0_translator_avalon_anti_slave_0_write;                                                 // wave_gen_2_s0_translator:av_write -> wave_gen_2:avs_s0_write
	wire          wave_gen_2_s0_translator_avalon_anti_slave_0_read;                                                  // wave_gen_2_s0_translator:av_read -> wave_gen_2:avs_s0_read
	wire   [31:0] wave_gen_2_s0_translator_avalon_anti_slave_0_readdata;                                              // wave_gen_2:avs_s0_readdata -> wave_gen_2_s0_translator:av_readdata
	wire    [0:0] cpu_ddr2_clock_bridge_m0_burstcount;                                                                // cpu_ddr2_clock_bridge:m0_burstcount -> cpu_ddr2_clock_bridge_m0_translator:av_burstcount
	wire          cpu_ddr2_clock_bridge_m0_waitrequest;                                                               // cpu_ddr2_clock_bridge_m0_translator:av_waitrequest -> cpu_ddr2_clock_bridge:m0_waitrequest
	wire   [25:0] cpu_ddr2_clock_bridge_m0_address;                                                                   // cpu_ddr2_clock_bridge:m0_address -> cpu_ddr2_clock_bridge_m0_translator:av_address
	wire   [31:0] cpu_ddr2_clock_bridge_m0_writedata;                                                                 // cpu_ddr2_clock_bridge:m0_writedata -> cpu_ddr2_clock_bridge_m0_translator:av_writedata
	wire          cpu_ddr2_clock_bridge_m0_write;                                                                     // cpu_ddr2_clock_bridge:m0_write -> cpu_ddr2_clock_bridge_m0_translator:av_write
	wire          cpu_ddr2_clock_bridge_m0_read;                                                                      // cpu_ddr2_clock_bridge:m0_read -> cpu_ddr2_clock_bridge_m0_translator:av_read
	wire   [31:0] cpu_ddr2_clock_bridge_m0_readdata;                                                                  // cpu_ddr2_clock_bridge_m0_translator:av_readdata -> cpu_ddr2_clock_bridge:m0_readdata
	wire          cpu_ddr2_clock_bridge_m0_debugaccess;                                                               // cpu_ddr2_clock_bridge:m0_debugaccess -> cpu_ddr2_clock_bridge_m0_translator:av_debugaccess
	wire    [3:0] cpu_ddr2_clock_bridge_m0_byteenable;                                                                // cpu_ddr2_clock_bridge:m0_byteenable -> cpu_ddr2_clock_bridge_m0_translator:av_byteenable
	wire          cpu_ddr2_clock_bridge_m0_readdatavalid;                                                             // cpu_ddr2_clock_bridge_m0_translator:av_readdatavalid -> cpu_ddr2_clock_bridge:m0_readdatavalid
	wire          ddr2_s1_translator_avalon_anti_slave_0_waitrequest;                                                 // ddr2:local_ready -> ddr2_s1_translator:av_waitrequest
	wire    [2:0] ddr2_s1_translator_avalon_anti_slave_0_burstcount;                                                  // ddr2_s1_translator:av_burstcount -> ddr2:local_size
	wire   [31:0] ddr2_s1_translator_avalon_anti_slave_0_writedata;                                                   // ddr2_s1_translator:av_writedata -> ddr2:local_wdata
	wire   [23:0] ddr2_s1_translator_avalon_anti_slave_0_address;                                                     // ddr2_s1_translator:av_address -> ddr2:local_address
	wire          ddr2_s1_translator_avalon_anti_slave_0_write;                                                       // ddr2_s1_translator:av_write -> ddr2:local_write_req
	wire          ddr2_s1_translator_avalon_anti_slave_0_beginbursttransfer;                                          // ddr2_s1_translator:av_beginbursttransfer -> ddr2:local_burstbegin
	wire          ddr2_s1_translator_avalon_anti_slave_0_read;                                                        // ddr2_s1_translator:av_read -> ddr2:local_read_req
	wire   [31:0] ddr2_s1_translator_avalon_anti_slave_0_readdata;                                                    // ddr2:local_rdata -> ddr2_s1_translator:av_readdata
	wire          ddr2_s1_translator_avalon_anti_slave_0_readdatavalid;                                               // ddr2:local_rdata_valid -> ddr2_s1_translator:av_readdatavalid
	wire    [3:0] ddr2_s1_translator_avalon_anti_slave_0_byteenable;                                                  // ddr2_s1_translator:av_byteenable -> ddr2:local_be
	wire          ddr2_reset_request_n_reset;                                                                         // ddr2:reset_request_n -> [ddr2_s1_translator:reset, ddr2_s1_translator_avalon_universal_slave_0_agent:reset, ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_030:reset, rsp_xbar_demux_030:reset, rst_controller:reset_in2, rst_controller_001:reset_in2, rst_controller_002:reset_in2, rst_controller_004:reset_in2, rst_controller_005:reset_in2]
	wire          nios2_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // nios2_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios2_instruction_master_translator_avalon_universal_master_0_burstcount;                           // nios2_instruction_master_translator:uav_burstcount -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_instruction_master_translator_avalon_universal_master_0_writedata;                            // nios2_instruction_master_translator:uav_writedata -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [26:0] nios2_instruction_master_translator_avalon_universal_master_0_address;                              // nios2_instruction_master_translator:uav_address -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_instruction_master_translator_avalon_universal_master_0_lock;                                 // nios2_instruction_master_translator:uav_lock -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_instruction_master_translator_avalon_universal_master_0_write;                                // nios2_instruction_master_translator:uav_write -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_instruction_master_translator_avalon_universal_master_0_read;                                 // nios2_instruction_master_translator:uav_read -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_instruction_master_translator_avalon_universal_master_0_readdata;                             // nios2_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_instruction_master_translator:uav_readdata
	wire          nios2_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // nios2_instruction_master_translator:uav_debugaccess -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_instruction_master_translator_avalon_universal_master_0_byteenable;                           // nios2_instruction_master_translator:uav_byteenable -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // nios2_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_instruction_master_translator:uav_readdatavalid
	wire          nios2_data_master_translator_avalon_universal_master_0_waitrequest;                                 // nios2_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_data_master_translator:uav_waitrequest
	wire    [2:0] nios2_data_master_translator_avalon_universal_master_0_burstcount;                                  // nios2_data_master_translator:uav_burstcount -> nios2_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_data_master_translator_avalon_universal_master_0_writedata;                                   // nios2_data_master_translator:uav_writedata -> nios2_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [26:0] nios2_data_master_translator_avalon_universal_master_0_address;                                     // nios2_data_master_translator:uav_address -> nios2_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_data_master_translator_avalon_universal_master_0_lock;                                        // nios2_data_master_translator:uav_lock -> nios2_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_data_master_translator_avalon_universal_master_0_write;                                       // nios2_data_master_translator:uav_write -> nios2_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_data_master_translator_avalon_universal_master_0_read;                                        // nios2_data_master_translator:uav_read -> nios2_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_data_master_translator_avalon_universal_master_0_readdata;                                    // nios2_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_data_master_translator:uav_readdata
	wire          nios2_data_master_translator_avalon_universal_master_0_debugaccess;                                 // nios2_data_master_translator:uav_debugaccess -> nios2_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_data_master_translator_avalon_universal_master_0_byteenable;                                  // nios2_data_master_translator:uav_byteenable -> nios2_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_data_master_translator_avalon_universal_master_0_readdatavalid;                               // nios2_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_data_master_translator:uav_readdatavalid
	wire          dma_0_read_master_translator_avalon_universal_master_0_waitrequest;                                 // dma_0_read_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_0_read_master_translator:uav_waitrequest
	wire    [2:0] dma_0_read_master_translator_avalon_universal_master_0_burstcount;                                  // dma_0_read_master_translator:uav_burstcount -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] dma_0_read_master_translator_avalon_universal_master_0_writedata;                                   // dma_0_read_master_translator:uav_writedata -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [26:0] dma_0_read_master_translator_avalon_universal_master_0_address;                                     // dma_0_read_master_translator:uav_address -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_0_read_master_translator_avalon_universal_master_0_lock;                                        // dma_0_read_master_translator:uav_lock -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_0_read_master_translator_avalon_universal_master_0_write;                                       // dma_0_read_master_translator:uav_write -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_0_read_master_translator_avalon_universal_master_0_read;                                        // dma_0_read_master_translator:uav_read -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] dma_0_read_master_translator_avalon_universal_master_0_readdata;                                    // dma_0_read_master_translator_avalon_universal_master_0_agent:av_readdata -> dma_0_read_master_translator:uav_readdata
	wire          dma_0_read_master_translator_avalon_universal_master_0_debugaccess;                                 // dma_0_read_master_translator:uav_debugaccess -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] dma_0_read_master_translator_avalon_universal_master_0_byteenable;                                  // dma_0_read_master_translator:uav_byteenable -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_0_read_master_translator_avalon_universal_master_0_readdatavalid;                               // dma_0_read_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_0_read_master_translator:uav_readdatavalid
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // nios2_jtag_debug_module_translator:uav_waitrequest -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_jtag_debug_module_translator:uav_writedata
	wire   [26:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_jtag_debug_module_translator:uav_address
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_jtag_debug_module_translator:uav_write
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_jtag_debug_module_translator:uav_lock
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // nios2_jtag_debug_module_translator:uav_readdata -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // nios2_jtag_debug_module_translator:uav_readdatavalid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_jtag_debug_module_translator:uav_byteenable
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [100:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [100:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // epcs_flash_epcs_control_port_translator:uav_waitrequest -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;               // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> epcs_flash_epcs_control_port_translator:uav_burstcount
	wire   [31:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;                // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> epcs_flash_epcs_control_port_translator:uav_writedata
	wire   [26:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address;                  // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_address -> epcs_flash_epcs_control_port_translator:uav_address
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write;                    // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_write -> epcs_flash_epcs_control_port_translator:uav_write
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                     // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> epcs_flash_epcs_control_port_translator:uav_lock
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read;                     // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_read -> epcs_flash_epcs_control_port_translator:uav_read
	wire   [31:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                 // epcs_flash_epcs_control_port_translator:uav_readdata -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // epcs_flash_epcs_control_port_translator:uav_readdatavalid -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> epcs_flash_epcs_control_port_translator:uav_debugaccess
	wire    [3:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;               // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> epcs_flash_epcs_control_port_translator:uav_byteenable
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;             // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [100:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;              // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;             // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [100:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // onchip_ram_s1_translator:uav_waitrequest -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_ram_s1_translator:uav_burstcount
	wire   [31:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_ram_s1_translator:uav_writedata
	wire   [26:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_ram_s1_translator:uav_address
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_ram_s1_translator:uav_write
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_ram_s1_translator:uav_lock
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_ram_s1_translator:uav_read
	wire   [31:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // onchip_ram_s1_translator:uav_readdata -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // onchip_ram_s1_translator:uav_readdatavalid -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_ram_s1_translator:uav_debugaccess
	wire    [3:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_ram_s1_translator:uav_byteenable
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [100:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [100:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // cpu_ddr2_clock_bridge_s0_translator:uav_waitrequest -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_ddr2_clock_bridge_s0_translator:uav_burstcount
	wire   [31:0] cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                    // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_ddr2_clock_bridge_s0_translator:uav_writedata
	wire   [26:0] cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                      // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> cpu_ddr2_clock_bridge_s0_translator:uav_address
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                        // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> cpu_ddr2_clock_bridge_s0_translator:uav_write
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                         // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_ddr2_clock_bridge_s0_translator:uav_lock
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                         // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> cpu_ddr2_clock_bridge_s0_translator:uav_read
	wire   [31:0] cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                     // cpu_ddr2_clock_bridge_s0_translator:uav_readdata -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // cpu_ddr2_clock_bridge_s0_translator:uav_readdatavalid -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_ddr2_clock_bridge_s0_translator:uav_debugaccess
	wire    [3:0] cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_ddr2_clock_bridge_s0_translator:uav_byteenable
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [100:0] cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                  // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [100:0] cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // slow_peripheral_bridge_s0_translator:uav_waitrequest -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> slow_peripheral_bridge_s0_translator:uav_burstcount
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                   // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> slow_peripheral_bridge_s0_translator:uav_writedata
	wire   [26:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                     // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> slow_peripheral_bridge_s0_translator:uav_address
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                       // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> slow_peripheral_bridge_s0_translator:uav_write
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                        // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> slow_peripheral_bridge_s0_translator:uav_lock
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                        // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> slow_peripheral_bridge_s0_translator:uav_read
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                    // slow_peripheral_bridge_s0_translator:uav_readdata -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // slow_peripheral_bridge_s0_translator:uav_readdatavalid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> slow_peripheral_bridge_s0_translator:uav_debugaccess
	wire    [3:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> slow_peripheral_bridge_s0_translator:uav_byteenable
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [100:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                 // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [100:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // dma_0_control_port_slave_translator:uav_waitrequest -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> dma_0_control_port_slave_translator:uav_burstcount
	wire   [31:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                    // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> dma_0_control_port_slave_translator:uav_writedata
	wire   [26:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                      // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> dma_0_control_port_slave_translator:uav_address
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                        // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> dma_0_control_port_slave_translator:uav_write
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                         // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> dma_0_control_port_slave_translator:uav_lock
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                         // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> dma_0_control_port_slave_translator:uav_read
	wire   [31:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                     // dma_0_control_port_slave_translator:uav_readdata -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // dma_0_control_port_slave_translator:uav_readdatavalid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dma_0_control_port_slave_translator:uav_debugaccess
	wire    [3:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> dma_0_control_port_slave_translator:uav_byteenable
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [100:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                  // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [100:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest;                         // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> slow_peripheral_bridge_m0_translator:uav_waitrequest
	wire    [2:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount;                          // slow_peripheral_bridge_m0_translator:uav_burstcount -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_writedata;                           // slow_peripheral_bridge_m0_translator:uav_writedata -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire    [9:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_address;                             // slow_peripheral_bridge_m0_translator:uav_address -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_lock;                                // slow_peripheral_bridge_m0_translator:uav_lock -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_write;                               // slow_peripheral_bridge_m0_translator:uav_write -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_read;                                // slow_peripheral_bridge_m0_translator:uav_read -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdata;                            // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> slow_peripheral_bridge_m0_translator:uav_readdata
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess;                         // slow_peripheral_bridge_m0_translator:uav_debugaccess -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable;                          // slow_peripheral_bridge_m0_translator:uav_byteenable -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                       // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> slow_peripheral_bridge_m0_translator:uav_readdatavalid
	wire          dma_0_write_master_translator_avalon_universal_master_0_waitrequest;                                // dma_0_write_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_0_write_master_translator:uav_waitrequest
	wire    [2:0] dma_0_write_master_translator_avalon_universal_master_0_burstcount;                                 // dma_0_write_master_translator:uav_burstcount -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] dma_0_write_master_translator_avalon_universal_master_0_writedata;                                  // dma_0_write_master_translator:uav_writedata -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_writedata
	wire    [9:0] dma_0_write_master_translator_avalon_universal_master_0_address;                                    // dma_0_write_master_translator:uav_address -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_0_write_master_translator_avalon_universal_master_0_lock;                                       // dma_0_write_master_translator:uav_lock -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_0_write_master_translator_avalon_universal_master_0_write;                                      // dma_0_write_master_translator:uav_write -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_0_write_master_translator_avalon_universal_master_0_read;                                       // dma_0_write_master_translator:uav_read -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] dma_0_write_master_translator_avalon_universal_master_0_readdata;                                   // dma_0_write_master_translator_avalon_universal_master_0_agent:av_readdata -> dma_0_write_master_translator:uav_readdata
	wire          dma_0_write_master_translator_avalon_universal_master_0_debugaccess;                                // dma_0_write_master_translator:uav_debugaccess -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] dma_0_write_master_translator_avalon_universal_master_0_byteenable;                                 // dma_0_write_master_translator:uav_byteenable -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_0_write_master_translator_avalon_universal_master_0_readdatavalid;                              // dma_0_write_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_0_write_master_translator:uav_readdatavalid
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // altpll_0_pll_slave_translator:uav_waitrequest -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> altpll_0_pll_slave_translator:uav_burstcount
	wire   [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> altpll_0_pll_slave_translator:uav_writedata
	wire    [9:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> altpll_0_pll_slave_translator:uav_address
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> altpll_0_pll_slave_translator:uav_write
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> altpll_0_pll_slave_translator:uav_lock
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> altpll_0_pll_slave_translator:uav_read
	wire   [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // altpll_0_pll_slave_translator:uav_readdata -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // altpll_0_pll_slave_translator:uav_readdatavalid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> altpll_0_pll_slave_translator:uav_debugaccess
	wire    [3:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> altpll_0_pll_slave_translator:uav_byteenable
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                  // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                   // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                  // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire    [9:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                          // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire    [9:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // systimer_s1_translator:uav_waitrequest -> systimer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] systimer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // systimer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> systimer_s1_translator:uav_burstcount
	wire   [31:0] systimer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // systimer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> systimer_s1_translator:uav_writedata
	wire    [9:0] systimer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // systimer_s1_translator_avalon_universal_slave_0_agent:m0_address -> systimer_s1_translator:uav_address
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // systimer_s1_translator_avalon_universal_slave_0_agent:m0_write -> systimer_s1_translator:uav_write
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // systimer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> systimer_s1_translator:uav_lock
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // systimer_s1_translator_avalon_universal_slave_0_agent:m0_read -> systimer_s1_translator:uav_read
	wire   [31:0] systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // systimer_s1_translator:uav_readdata -> systimer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // systimer_s1_translator:uav_readdatavalid -> systimer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // systimer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> systimer_s1_translator:uav_debugaccess
	wire    [3:0] systimer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // systimer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> systimer_s1_translator:uav_byteenable
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // systimer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // systimer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // systimer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // systimer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> systimer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> systimer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> systimer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // systimer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                         // systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                          // systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                         // systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // pio_key_s1_translator:uav_waitrequest -> pio_key_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_key_s1_translator:uav_burstcount
	wire   [31:0] pio_key_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_key_s1_translator:uav_writedata
	wire    [9:0] pio_key_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_key_s1_translator:uav_address
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_key_s1_translator:uav_write
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_key_s1_translator:uav_lock
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_key_s1_translator:uav_read
	wire   [31:0] pio_key_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // pio_key_s1_translator:uav_readdata -> pio_key_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // pio_key_s1_translator:uav_readdatavalid -> pio_key_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_key_s1_translator:uav_debugaccess
	wire    [3:0] pio_key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_key_s1_translator:uav_byteenable
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // pio_key_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // pio_key_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // pio_key_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // pio_key_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_key_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_key_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_key_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_key_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_key_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // pio_key_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // pio_key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // pio_key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> pio_key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                          // pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> pio_key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                           // pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> pio_key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                          // pio_key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // spi_0_spi_control_port_translator:uav_waitrequest -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> spi_0_spi_control_port_translator:uav_burstcount
	wire   [31:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;                      // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> spi_0_spi_control_port_translator:uav_writedata
	wire    [9:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address;                        // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_address -> spi_0_spi_control_port_translator:uav_address
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write;                          // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_write -> spi_0_spi_control_port_translator:uav_write
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                           // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> spi_0_spi_control_port_translator:uav_lock
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read;                           // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_read -> spi_0_spi_control_port_translator:uav_read
	wire   [31:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                       // spi_0_spi_control_port_translator:uav_readdata -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // spi_0_spi_control_port_translator:uav_readdatavalid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> spi_0_spi_control_port_translator:uav_debugaccess
	wire    [3:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> spi_0_spi_control_port_translator:uav_byteenable
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;                    // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;              // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;               // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;              // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // uart_0_s1_translator:uav_waitrequest -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart_0_s1_translator:uav_burstcount
	wire   [31:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart_0_s1_translator:uav_writedata
	wire    [9:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart_0_s1_translator:uav_address
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart_0_s1_translator:uav_write
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart_0_s1_translator:uav_lock
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart_0_s1_translator:uav_read
	wire   [31:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // uart_0_s1_translator:uav_readdata -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // uart_0_s1_translator:uav_readdatavalid -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart_0_s1_translator:uav_debugaccess
	wire    [3:0] uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // uart_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart_0_s1_translator:uav_byteenable
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                           // uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                            // uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                           // uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // pio_led_s1_translator:uav_waitrequest -> pio_led_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_led_s1_translator:uav_burstcount
	wire   [31:0] pio_led_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_led_s1_translator:uav_writedata
	wire    [9:0] pio_led_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_led_s1_translator:uav_address
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_led_s1_translator:uav_write
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_led_s1_translator:uav_lock
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_led_s1_translator:uav_read
	wire   [31:0] pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // pio_led_s1_translator:uav_readdata -> pio_led_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // pio_led_s1_translator:uav_readdatavalid -> pio_led_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_led_s1_translator:uav_debugaccess
	wire    [3:0] pio_led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_led_s1_translator:uav_byteenable
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // pio_led_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // pio_led_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // pio_led_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // pio_led_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_led_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // pio_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                          // pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                           // pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                          // pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // timestamp_s1_translator:uav_waitrequest -> timestamp_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timestamp_s1_translator:uav_burstcount
	wire   [31:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timestamp_s1_translator:uav_writedata
	wire    [9:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_address -> timestamp_s1_translator:uav_address
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_write -> timestamp_s1_translator:uav_write
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timestamp_s1_translator:uav_lock
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_read -> timestamp_s1_translator:uav_read
	wire   [31:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // timestamp_s1_translator:uav_readdata -> timestamp_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // timestamp_s1_translator:uav_readdatavalid -> timestamp_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timestamp_s1_translator:uav_debugaccess
	wire    [3:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timestamp_s1_translator:uav_byteenable
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                        // timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                         // timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                        // timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // spi_ad5781_spi_control_port_translator:uav_waitrequest -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;                // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> spi_ad5781_spi_control_port_translator:uav_burstcount
	wire   [31:0] spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;                 // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> spi_ad5781_spi_control_port_translator:uav_writedata
	wire    [9:0] spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address;                   // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:m0_address -> spi_ad5781_spi_control_port_translator:uav_address
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write;                     // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:m0_write -> spi_ad5781_spi_control_port_translator:uav_write
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                      // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> spi_ad5781_spi_control_port_translator:uav_lock
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read;                      // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:m0_read -> spi_ad5781_spi_control_port_translator:uav_read
	wire   [31:0] spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                  // spi_ad5781_spi_control_port_translator:uav_readdata -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // spi_ad5781_spi_control_port_translator:uav_readdatavalid -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> spi_ad5781_spi_control_port_translator:uav_debugaccess
	wire    [3:0] spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;                // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> spi_ad5781_spi_control_port_translator:uav_byteenable
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;              // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;               // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;              // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;         // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;          // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;         // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // ad9245_2_s1_translator:uav_waitrequest -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // ad9245_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ad9245_2_s1_translator:uav_burstcount
	wire   [31:0] ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // ad9245_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ad9245_2_s1_translator:uav_writedata
	wire    [9:0] ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // ad9245_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> ad9245_2_s1_translator:uav_address
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // ad9245_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> ad9245_2_s1_translator:uav_write
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // ad9245_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ad9245_2_s1_translator:uav_lock
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // ad9245_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> ad9245_2_s1_translator:uav_read
	wire   [31:0] ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // ad9245_2_s1_translator:uav_readdata -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // ad9245_2_s1_translator:uav_readdatavalid -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // ad9245_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ad9245_2_s1_translator:uav_debugaccess
	wire    [3:0] ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // ad9245_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ad9245_2_s1_translator:uav_byteenable
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // ad9245_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // ad9245_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // ad9245_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] ad9245_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // ad9245_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // ad9245_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // ad9245_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // ad9245_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                         // ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                          // ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                         // ad9245_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // clk_gen_s1_translator:uav_waitrequest -> clk_gen_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // clk_gen_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> clk_gen_s1_translator:uav_burstcount
	wire   [31:0] clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // clk_gen_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> clk_gen_s1_translator:uav_writedata
	wire    [9:0] clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // clk_gen_s1_translator_avalon_universal_slave_0_agent:m0_address -> clk_gen_s1_translator:uav_address
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // clk_gen_s1_translator_avalon_universal_slave_0_agent:m0_write -> clk_gen_s1_translator:uav_write
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // clk_gen_s1_translator_avalon_universal_slave_0_agent:m0_lock -> clk_gen_s1_translator:uav_lock
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // clk_gen_s1_translator_avalon_universal_slave_0_agent:m0_read -> clk_gen_s1_translator:uav_read
	wire   [31:0] clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // clk_gen_s1_translator:uav_readdata -> clk_gen_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // clk_gen_s1_translator:uav_readdatavalid -> clk_gen_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // clk_gen_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> clk_gen_s1_translator:uav_debugaccess
	wire    [3:0] clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // clk_gen_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> clk_gen_s1_translator:uav_byteenable
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // clk_gen_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // clk_gen_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // clk_gen_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] clk_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // clk_gen_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> clk_gen_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> clk_gen_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> clk_gen_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> clk_gen_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> clk_gen_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // clk_gen_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // clk_gen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // clk_gen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> clk_gen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                          // clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> clk_gen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                           // clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> clk_gen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                          // clk_gen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // oc_i2c_master_0_s1_translator:uav_waitrequest -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> oc_i2c_master_0_s1_translator:uav_burstcount
	wire   [31:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> oc_i2c_master_0_s1_translator:uav_writedata
	wire    [9:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> oc_i2c_master_0_s1_translator:uav_address
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> oc_i2c_master_0_s1_translator:uav_write
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> oc_i2c_master_0_s1_translator:uav_lock
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> oc_i2c_master_0_s1_translator:uav_read
	wire   [31:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // oc_i2c_master_0_s1_translator:uav_readdata -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // oc_i2c_master_0_s1_translator:uav_readdatavalid -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> oc_i2c_master_0_s1_translator:uav_debugaccess
	wire    [3:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> oc_i2c_master_0_s1_translator:uav_byteenable
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                  // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                   // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                  // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // spi_master_0_s1_translator:uav_waitrequest -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // spi_master_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> spi_master_0_s1_translator:uav_burstcount
	wire   [31:0] spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // spi_master_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> spi_master_0_s1_translator:uav_writedata
	wire    [9:0] spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // spi_master_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> spi_master_0_s1_translator:uav_address
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // spi_master_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> spi_master_0_s1_translator:uav_write
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // spi_master_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> spi_master_0_s1_translator:uav_lock
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // spi_master_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> spi_master_0_s1_translator:uav_read
	wire   [31:0] spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // spi_master_0_s1_translator:uav_readdata -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // spi_master_0_s1_translator:uav_readdatavalid -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // spi_master_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> spi_master_0_s1_translator:uav_debugaccess
	wire    [3:0] spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // spi_master_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> spi_master_0_s1_translator:uav_byteenable
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // spi_master_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // spi_master_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // spi_master_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] spi_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // spi_master_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // spi_master_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // spi_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // spi_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                     // spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                      // spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                     // spi_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // ad9266_spi_control_port_translator:uav_waitrequest -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> ad9266_spi_control_port_translator:uav_burstcount
	wire   [31:0] ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;                     // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> ad9266_spi_control_port_translator:uav_writedata
	wire    [9:0] ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address;                       // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:m0_address -> ad9266_spi_control_port_translator:uav_address
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write;                         // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:m0_write -> ad9266_spi_control_port_translator:uav_write
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                          // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> ad9266_spi_control_port_translator:uav_lock
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read;                          // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:m0_read -> ad9266_spi_control_port_translator:uav_read
	wire   [31:0] ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                      // ad9266_spi_control_port_translator:uav_readdata -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // ad9266_spi_control_port_translator:uav_readdatavalid -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ad9266_spi_control_port_translator:uav_debugaccess
	wire    [3:0] ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> ad9266_spi_control_port_translator:uav_byteenable
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;                   // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;             // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;              // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;             // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // ad9245_1_s1_translator:uav_waitrequest -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // ad9245_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ad9245_1_s1_translator:uav_burstcount
	wire   [31:0] ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // ad9245_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ad9245_1_s1_translator:uav_writedata
	wire    [9:0] ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // ad9245_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> ad9245_1_s1_translator:uav_address
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // ad9245_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> ad9245_1_s1_translator:uav_write
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // ad9245_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ad9245_1_s1_translator:uav_lock
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // ad9245_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> ad9245_1_s1_translator:uav_read
	wire   [31:0] ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // ad9245_1_s1_translator:uav_readdata -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // ad9245_1_s1_translator:uav_readdatavalid -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // ad9245_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ad9245_1_s1_translator:uav_debugaccess
	wire    [3:0] ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // ad9245_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ad9245_1_s1_translator:uav_byteenable
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // ad9245_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // ad9245_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // ad9245_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] ad9245_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // ad9245_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // ad9245_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // ad9245_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // ad9245_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                         // ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                          // ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                         // ad9245_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // dac2904_1_s0_translator:uav_waitrequest -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // dac2904_1_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> dac2904_1_s0_translator:uav_burstcount
	wire   [31:0] dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                                // dac2904_1_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> dac2904_1_s0_translator:uav_writedata
	wire    [9:0] dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_address;                                  // dac2904_1_s0_translator_avalon_universal_slave_0_agent:m0_address -> dac2904_1_s0_translator:uav_address
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_write;                                    // dac2904_1_s0_translator_avalon_universal_slave_0_agent:m0_write -> dac2904_1_s0_translator:uav_write
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                     // dac2904_1_s0_translator_avalon_universal_slave_0_agent:m0_lock -> dac2904_1_s0_translator:uav_lock
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_read;                                     // dac2904_1_s0_translator_avalon_universal_slave_0_agent:m0_read -> dac2904_1_s0_translator:uav_read
	wire   [31:0] dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // dac2904_1_s0_translator:uav_readdata -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // dac2904_1_s0_translator:uav_readdatavalid -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // dac2904_1_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dac2904_1_s0_translator:uav_debugaccess
	wire    [3:0] dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // dac2904_1_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> dac2904_1_s0_translator:uav_byteenable
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // dac2904_1_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // dac2904_1_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // dac2904_1_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] dac2904_1_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                              // dac2904_1_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // dac2904_1_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // dac2904_1_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // dac2904_1_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                        // dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                         // dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                        // dac2904_1_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // dac2904_2_s0_translator:uav_waitrequest -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // dac2904_2_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> dac2904_2_s0_translator:uav_burstcount
	wire   [31:0] dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                                // dac2904_2_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> dac2904_2_s0_translator:uav_writedata
	wire    [9:0] dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_address;                                  // dac2904_2_s0_translator_avalon_universal_slave_0_agent:m0_address -> dac2904_2_s0_translator:uav_address
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_write;                                    // dac2904_2_s0_translator_avalon_universal_slave_0_agent:m0_write -> dac2904_2_s0_translator:uav_write
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                     // dac2904_2_s0_translator_avalon_universal_slave_0_agent:m0_lock -> dac2904_2_s0_translator:uav_lock
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_read;                                     // dac2904_2_s0_translator_avalon_universal_slave_0_agent:m0_read -> dac2904_2_s0_translator:uav_read
	wire   [31:0] dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // dac2904_2_s0_translator:uav_readdata -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // dac2904_2_s0_translator:uav_readdatavalid -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // dac2904_2_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dac2904_2_s0_translator:uav_debugaccess
	wire    [3:0] dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // dac2904_2_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> dac2904_2_s0_translator:uav_byteenable
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // dac2904_2_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // dac2904_2_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // dac2904_2_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] dac2904_2_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                              // dac2904_2_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // dac2904_2_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // dac2904_2_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // dac2904_2_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                        // dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                         // dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                        // dac2904_2_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // dac2904_3_s0_translator:uav_waitrequest -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // dac2904_3_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> dac2904_3_s0_translator:uav_burstcount
	wire   [31:0] dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                                // dac2904_3_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> dac2904_3_s0_translator:uav_writedata
	wire    [9:0] dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_address;                                  // dac2904_3_s0_translator_avalon_universal_slave_0_agent:m0_address -> dac2904_3_s0_translator:uav_address
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_write;                                    // dac2904_3_s0_translator_avalon_universal_slave_0_agent:m0_write -> dac2904_3_s0_translator:uav_write
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                     // dac2904_3_s0_translator_avalon_universal_slave_0_agent:m0_lock -> dac2904_3_s0_translator:uav_lock
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_read;                                     // dac2904_3_s0_translator_avalon_universal_slave_0_agent:m0_read -> dac2904_3_s0_translator:uav_read
	wire   [31:0] dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // dac2904_3_s0_translator:uav_readdata -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // dac2904_3_s0_translator:uav_readdatavalid -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // dac2904_3_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dac2904_3_s0_translator:uav_debugaccess
	wire    [3:0] dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // dac2904_3_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> dac2904_3_s0_translator:uav_byteenable
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // dac2904_3_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // dac2904_3_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // dac2904_3_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] dac2904_3_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                              // dac2904_3_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // dac2904_3_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // dac2904_3_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // dac2904_3_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                        // dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                         // dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                        // dac2904_3_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // dac2904_4_s0_translator:uav_waitrequest -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // dac2904_4_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> dac2904_4_s0_translator:uav_burstcount
	wire   [31:0] dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                                // dac2904_4_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> dac2904_4_s0_translator:uav_writedata
	wire    [9:0] dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_address;                                  // dac2904_4_s0_translator_avalon_universal_slave_0_agent:m0_address -> dac2904_4_s0_translator:uav_address
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_write;                                    // dac2904_4_s0_translator_avalon_universal_slave_0_agent:m0_write -> dac2904_4_s0_translator:uav_write
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                     // dac2904_4_s0_translator_avalon_universal_slave_0_agent:m0_lock -> dac2904_4_s0_translator:uav_lock
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_read;                                     // dac2904_4_s0_translator_avalon_universal_slave_0_agent:m0_read -> dac2904_4_s0_translator:uav_read
	wire   [31:0] dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // dac2904_4_s0_translator:uav_readdata -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // dac2904_4_s0_translator:uav_readdatavalid -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // dac2904_4_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dac2904_4_s0_translator:uav_debugaccess
	wire    [3:0] dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // dac2904_4_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> dac2904_4_s0_translator:uav_byteenable
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // dac2904_4_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // dac2904_4_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // dac2904_4_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] dac2904_4_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                              // dac2904_4_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // dac2904_4_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // dac2904_4_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // dac2904_4_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                        // dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                         // dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                        // dac2904_4_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // wave_gen_0_s0_translator:uav_waitrequest -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> wave_gen_0_s0_translator:uav_burstcount
	wire   [31:0] wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                               // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> wave_gen_0_s0_translator:uav_writedata
	wire    [9:0] wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_address;                                 // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:m0_address -> wave_gen_0_s0_translator:uav_address
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_write;                                   // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:m0_write -> wave_gen_0_s0_translator:uav_write
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                    // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:m0_lock -> wave_gen_0_s0_translator:uav_lock
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_read;                                    // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:m0_read -> wave_gen_0_s0_translator:uav_read
	wire   [31:0] wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                // wave_gen_0_s0_translator:uav_readdata -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // wave_gen_0_s0_translator:uav_readdatavalid -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> wave_gen_0_s0_translator:uav_debugaccess
	wire    [3:0] wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> wave_gen_0_s0_translator:uav_byteenable
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                             // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                       // wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                        // wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                       // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // demodulation_0_s0_translator:uav_waitrequest -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // demodulation_0_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> demodulation_0_s0_translator:uav_burstcount
	wire   [31:0] demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                           // demodulation_0_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> demodulation_0_s0_translator:uav_writedata
	wire    [9:0] demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_address;                             // demodulation_0_s0_translator_avalon_universal_slave_0_agent:m0_address -> demodulation_0_s0_translator:uav_address
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_write;                               // demodulation_0_s0_translator_avalon_universal_slave_0_agent:m0_write -> demodulation_0_s0_translator:uav_write
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                // demodulation_0_s0_translator_avalon_universal_slave_0_agent:m0_lock -> demodulation_0_s0_translator:uav_lock
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_read;                                // demodulation_0_s0_translator_avalon_universal_slave_0_agent:m0_read -> demodulation_0_s0_translator:uav_read
	wire   [31:0] demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                            // demodulation_0_s0_translator:uav_readdata -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // demodulation_0_s0_translator:uav_readdatavalid -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // demodulation_0_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> demodulation_0_s0_translator:uav_debugaccess
	wire    [3:0] demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // demodulation_0_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> demodulation_0_s0_translator:uav_byteenable
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // demodulation_0_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // demodulation_0_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // demodulation_0_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] demodulation_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                         // demodulation_0_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // demodulation_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // demodulation_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // demodulation_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                   // demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                    // demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                   // demodulation_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // wave_gen_1_s0_translator:uav_waitrequest -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> wave_gen_1_s0_translator:uav_burstcount
	wire   [31:0] wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                               // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> wave_gen_1_s0_translator:uav_writedata
	wire    [9:0] wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_address;                                 // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:m0_address -> wave_gen_1_s0_translator:uav_address
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_write;                                   // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:m0_write -> wave_gen_1_s0_translator:uav_write
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                    // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:m0_lock -> wave_gen_1_s0_translator:uav_lock
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_read;                                    // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:m0_read -> wave_gen_1_s0_translator:uav_read
	wire   [31:0] wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                // wave_gen_1_s0_translator:uav_readdata -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // wave_gen_1_s0_translator:uav_readdatavalid -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> wave_gen_1_s0_translator:uav_debugaccess
	wire    [3:0] wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> wave_gen_1_s0_translator:uav_byteenable
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                             // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                       // wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                        // wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                       // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // wave_gen_2_s0_translator:uav_waitrequest -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> wave_gen_2_s0_translator:uav_burstcount
	wire   [31:0] wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                               // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> wave_gen_2_s0_translator:uav_writedata
	wire    [9:0] wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_address;                                 // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:m0_address -> wave_gen_2_s0_translator:uav_address
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_write;                                   // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:m0_write -> wave_gen_2_s0_translator:uav_write
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                    // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:m0_lock -> wave_gen_2_s0_translator:uav_lock
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_read;                                    // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:m0_read -> wave_gen_2_s0_translator:uav_read
	wire   [31:0] wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                                // wave_gen_2_s0_translator:uav_readdata -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // wave_gen_2_s0_translator:uav_readdatavalid -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> wave_gen_2_s0_translator:uav_debugaccess
	wire    [3:0] wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> wave_gen_2_s0_translator:uav_byteenable
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                             // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                       // wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                        // wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                       // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest;                          // cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_ddr2_clock_bridge_m0_translator:uav_waitrequest
	wire    [2:0] cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_burstcount;                           // cpu_ddr2_clock_bridge_m0_translator:uav_burstcount -> cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_writedata;                            // cpu_ddr2_clock_bridge_m0_translator:uav_writedata -> cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [25:0] cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_address;                              // cpu_ddr2_clock_bridge_m0_translator:uav_address -> cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_lock;                                 // cpu_ddr2_clock_bridge_m0_translator:uav_lock -> cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_write;                                // cpu_ddr2_clock_bridge_m0_translator:uav_write -> cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_read;                                 // cpu_ddr2_clock_bridge_m0_translator:uav_read -> cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_readdata;                             // cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> cpu_ddr2_clock_bridge_m0_translator:uav_readdata
	wire          cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess;                          // cpu_ddr2_clock_bridge_m0_translator:uav_debugaccess -> cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_byteenable;                           // cpu_ddr2_clock_bridge_m0_translator:uav_byteenable -> cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                        // cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_ddr2_clock_bridge_m0_translator:uav_readdatavalid
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // ddr2_s1_translator:uav_waitrequest -> ddr2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [4:0] ddr2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // ddr2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ddr2_s1_translator:uav_burstcount
	wire   [31:0] ddr2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // ddr2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ddr2_s1_translator:uav_writedata
	wire   [25:0] ddr2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // ddr2_s1_translator_avalon_universal_slave_0_agent:m0_address -> ddr2_s1_translator:uav_address
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // ddr2_s1_translator_avalon_universal_slave_0_agent:m0_write -> ddr2_s1_translator:uav_write
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // ddr2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ddr2_s1_translator:uav_lock
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // ddr2_s1_translator_avalon_universal_slave_0_agent:m0_read -> ddr2_s1_translator:uav_read
	wire   [31:0] ddr2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // ddr2_s1_translator:uav_readdata -> ddr2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // ddr2_s1_translator:uav_readdatavalid -> ddr2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // ddr2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ddr2_s1_translator:uav_debugaccess
	wire    [3:0] ddr2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // ddr2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ddr2_s1_translator:uav_byteenable
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // ddr2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // ddr2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // ddr2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [95:0] ddr2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // ddr2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ddr2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ddr2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ddr2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ddr2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [95:0] ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ddr2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // ddr2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // ddr2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ddr2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ddr2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // ddr2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ddr2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // ddr2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ddr2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire   [99:0] nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router:sink_ready -> nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // nios2_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          nios2_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // nios2_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          nios2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // nios2_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire   [99:0] nios2_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // nios2_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          nios2_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_001:sink_ready -> nios2_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          dma_0_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // dma_0_read_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          dma_0_read_master_translator_avalon_universal_master_0_agent_cp_valid;                              // dma_0_read_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          dma_0_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // dma_0_read_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire   [99:0] dma_0_read_master_translator_avalon_universal_master_0_agent_cp_data;                               // dma_0_read_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          dma_0_read_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_002:sink_ready -> dma_0_read_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire   [99:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router:sink_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                    // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [99:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data;                     // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_001:sink_ready -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire   [99:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_002:sink_ready -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                        // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire   [99:0] cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                         // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                        // id_router_003:sink_ready -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                       // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire   [99:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                        // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_004:sink_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                        // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire   [99:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                         // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                        // id_router_005:sink_ready -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                      // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;              // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire   [84:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                       // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                      // addr_router_003:sink_ready -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          dma_0_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // dma_0_write_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          dma_0_write_master_translator_avalon_universal_master_0_agent_cp_valid;                             // dma_0_write_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          dma_0_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // dma_0_write_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire   [84:0] dma_0_write_master_translator_avalon_universal_master_0_agent_cp_data;                              // dma_0_write_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          dma_0_write_master_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router_004:sink_ready -> dma_0_write_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire   [84:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_006:sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire   [84:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_007:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire   [84:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_008:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // systimer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // systimer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // systimer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire   [84:0] systimer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // systimer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_009:sink_ready -> systimer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // pio_key_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // pio_key_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // pio_key_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire   [84:0] pio_key_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // pio_key_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_010:sink_ready -> pio_key_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                          // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire   [84:0] spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data;                           // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_011:sink_ready -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire   [84:0] uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // uart_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_012:sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // pio_led_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // pio_led_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // pio_led_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire   [84:0] pio_led_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // pio_led_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_013:sink_ready -> pio_led_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire   [84:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_014:sink_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                     // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire   [84:0] spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data;                      // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                     // id_router_015:sink_ready -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // ad9245_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // ad9245_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // ad9245_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire   [84:0] ad9245_2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // ad9245_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          ad9245_2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_016:sink_ready -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // clk_gen_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // clk_gen_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // clk_gen_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire   [84:0] clk_gen_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // clk_gen_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          clk_gen_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_017:sink_ready -> clk_gen_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire   [84:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_018:sink_ready -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // spi_master_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // spi_master_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // spi_master_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire   [84:0] spi_master_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // spi_master_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire          spi_master_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_019:sink_ready -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                         // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire   [84:0] ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data;                          // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire          ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_020:sink_ready -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // ad9245_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // ad9245_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // ad9245_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire   [84:0] ad9245_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // ad9245_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire          ad9245_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_021:sink_ready -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // dac2904_1_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                    // dac2904_1_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // dac2904_1_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	wire   [84:0] dac2904_1_s0_translator_avalon_universal_slave_0_agent_rp_data;                                     // dac2904_1_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	wire          dac2904_1_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_022:sink_ready -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // dac2904_2_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_023:sink_endofpacket
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                    // dac2904_2_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_023:sink_valid
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // dac2904_2_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_023:sink_startofpacket
	wire   [84:0] dac2904_2_s0_translator_avalon_universal_slave_0_agent_rp_data;                                     // dac2904_2_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_023:sink_data
	wire          dac2904_2_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_023:sink_ready -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // dac2904_3_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_024:sink_endofpacket
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                    // dac2904_3_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_024:sink_valid
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // dac2904_3_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_024:sink_startofpacket
	wire   [84:0] dac2904_3_s0_translator_avalon_universal_slave_0_agent_rp_data;                                     // dac2904_3_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_024:sink_data
	wire          dac2904_3_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_024:sink_ready -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // dac2904_4_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_025:sink_endofpacket
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                    // dac2904_4_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_025:sink_valid
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // dac2904_4_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_025:sink_startofpacket
	wire   [84:0] dac2904_4_s0_translator_avalon_universal_slave_0_agent_rp_data;                                     // dac2904_4_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_025:sink_data
	wire          dac2904_4_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_025:sink_ready -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_026:sink_endofpacket
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                   // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_026:sink_valid
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_026:sink_startofpacket
	wire   [84:0] wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rp_data;                                    // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_026:sink_data
	wire          wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_026:sink_ready -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // demodulation_0_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_027:sink_endofpacket
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rp_valid;                               // demodulation_0_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_027:sink_valid
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // demodulation_0_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_027:sink_startofpacket
	wire   [84:0] demodulation_0_s0_translator_avalon_universal_slave_0_agent_rp_data;                                // demodulation_0_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_027:sink_data
	wire          demodulation_0_s0_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_027:sink_ready -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_028:sink_endofpacket
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                   // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_028:sink_valid
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_028:sink_startofpacket
	wire   [84:0] wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rp_data;                                    // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_028:sink_data
	wire          wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_028:sink_ready -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_029:sink_endofpacket
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                   // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_029:sink_valid
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_029:sink_startofpacket
	wire   [84:0] wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rp_data;                                    // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_029:sink_data
	wire          wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_029:sink_ready -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire          cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire          cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire   [94:0] cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire          cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_005:sink_ready -> cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // ddr2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_030:sink_endofpacket
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // ddr2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_030:sink_valid
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // ddr2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_030:sink_startofpacket
	wire   [94:0] ddr2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // ddr2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_030:sink_data
	wire          ddr2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_030:sink_ready -> ddr2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                        // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                              // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                      // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire   [99:0] addr_router_src_data;                                                                               // addr_router:src_data -> limiter:cmd_sink_data
	wire    [5:0] addr_router_src_channel;                                                                            // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                              // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                        // limiter:rsp_src_endofpacket -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                              // limiter:rsp_src_valid -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                      // limiter:rsp_src_startofpacket -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [99:0] limiter_rsp_src_data;                                                                               // limiter:rsp_src_data -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] limiter_rsp_src_channel;                                                                            // limiter:rsp_src_channel -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                              // nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_003_src_endofpacket;                                                                    // addr_router_003:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_003_src_valid;                                                                          // addr_router_003:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_003_src_startofpacket;                                                                  // addr_router_003:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire   [84:0] addr_router_003_src_data;                                                                           // addr_router_003:src_data -> limiter_001:cmd_sink_data
	wire   [23:0] addr_router_003_src_channel;                                                                        // addr_router_003:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_003_src_ready;                                                                          // limiter_001:cmd_sink_ready -> addr_router_003:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                    // limiter_001:rsp_src_endofpacket -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                          // limiter_001:rsp_src_valid -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                  // limiter_001:rsp_src_startofpacket -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [84:0] limiter_001_rsp_src_data;                                                                           // limiter_001:rsp_src_data -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire   [23:0] limiter_001_rsp_src_channel;                                                                        // limiter_001:rsp_src_channel -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                          // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          rst_controller_reset_out_reset;                                                                     // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_004:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_004:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cpu_ddr2_clock_bridge:s0_reset, cpu_ddr2_clock_bridge_s0_translator:reset, cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:reset, cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser_001:in_reset, crosser_002:in_reset, crosser_004:out_reset, crosser_005:out_reset, dma_0:system_reset_n, dma_0_control_port_slave_translator:reset, dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:reset, dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dma_0_read_master_translator:reset, dma_0_read_master_translator_avalon_universal_master_0_agent:reset, dma_0_write_master_translator:reset, dma_0_write_master_translator_avalon_universal_master_0_agent:reset, epcs_flash:reset_n, epcs_flash_epcs_control_port_translator:reset, epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:reset, epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, irq_synchronizer_005:sender_reset, irq_synchronizer_006:sender_reset, irq_synchronizer_007:sender_reset, irq_synchronizer_008:sender_reset, irq_synchronizer_009:sender_reset, limiter:reset, nios2:reset_n, nios2_data_master_translator:reset, nios2_data_master_translator_avalon_universal_master_0_agent:reset, nios2_instruction_master_translator:reset, nios2_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_jtag_debug_module_translator:reset, nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_ram:reset, onchip_ram_s1_translator:reset, onchip_ram_s1_translator_avalon_universal_slave_0_agent:reset, onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_004:reset, slow_peripheral_bridge:s0_reset, slow_peripheral_bridge_s0_translator:reset, slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:reset, slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          nios2_jtag_debug_module_reset_reset;                                                                // nios2:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_004:reset_in1, rst_controller_005:reset_in1]
	wire          rst_controller_001_reset_out_reset;                                                                 // rst_controller_001:reset_out -> [ad9245_1:reset_n, ad9245_1_s1_translator:reset, ad9245_1_s1_translator_avalon_universal_slave_0_agent:reset, ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ad9245_2:reset_n, ad9245_2_s1_translator:reset, ad9245_2_s1_translator_avalon_universal_slave_0_agent:reset, ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ad9266:reset_n, ad9266_spi_control_port_translator:reset, ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:reset, ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router_003:reset, clk_gen:reset_n, clk_gen_s1_translator:reset, clk_gen_s1_translator_avalon_universal_slave_0_agent:reset, clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux_003:reset, cmd_xbar_mux_021:reset, cmd_xbar_mux_022:reset, crosser:in_reset, crosser_001:out_reset, crosser_002:out_reset, crosser_003:out_reset, crosser_004:in_reset, crosser_005:in_reset, dac2904_1:reset_n, dac2904_1_s0_translator:reset, dac2904_1_s0_translator_avalon_universal_slave_0_agent:reset, dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dac2904_2:reset_n, dac2904_2_s0_translator:reset, dac2904_2_s0_translator_avalon_universal_slave_0_agent:reset, dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dac2904_3:reset_n, dac2904_3_s0_translator:reset, dac2904_3_s0_translator_avalon_universal_slave_0_agent:reset, dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dac2904_4:reset_n, dac2904_4_s0_translator:reset, dac2904_4_s0_translator_avalon_universal_slave_0_agent:reset, dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, demodulation_0:reset_n, demodulation_0_s0_translator:reset, demodulation_0_s0_translator_avalon_universal_slave_0_agent:reset, demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, id_router_022:reset, id_router_023:reset, id_router_024:reset, id_router_025:reset, id_router_026:reset, id_router_027:reset, id_router_028:reset, id_router_029:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, irq_synchronizer_005:receiver_reset, irq_synchronizer_006:receiver_reset, irq_synchronizer_007:receiver_reset, irq_synchronizer_008:receiver_reset, irq_synchronizer_009:receiver_reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter_001:reset, oc_i2c_master_0:wb_rst_i, oc_i2c_master_0_s1_translator:reset, oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:reset, oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_key:reset_n, pio_key_s1_translator:reset, pio_key_s1_translator_avalon_universal_slave_0_agent:reset, pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_led:reset_n, pio_led_s1_translator:reset, pio_led_s1_translator_avalon_universal_slave_0_agent:reset, pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_022:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_024:reset, rsp_xbar_demux_025:reset, rsp_xbar_demux_026:reset, rsp_xbar_demux_027:reset, rsp_xbar_demux_028:reset, rsp_xbar_demux_029:reset, rsp_xbar_mux_003:reset, slow_peripheral_bridge:m0_reset, slow_peripheral_bridge_m0_translator:reset, slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:reset, spi_0:reset_n, spi_0_spi_control_port_translator:reset, spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:reset, spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, spi_ad5781:reset_n, spi_ad5781_spi_control_port_translator:reset, spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:reset, spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, spi_master_0:reset_n, spi_master_0_s1_translator:reset, spi_master_0_s1_translator_avalon_universal_slave_0_agent:reset, spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, systimer:reset_n, systimer_s1_translator:reset, systimer_s1_translator_avalon_universal_slave_0_agent:reset, systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timestamp:reset_n, timestamp_s1_translator:reset, timestamp_s1_translator_avalon_universal_slave_0_agent:reset, timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, uart_0:reset_n, uart_0_s1_translator:reset, uart_0_s1_translator_avalon_universal_slave_0_agent:reset, uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, wave_gen_0:reset_n, wave_gen_0_s0_translator:reset, wave_gen_0_s0_translator_avalon_universal_slave_0_agent:reset, wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, wave_gen_1:reset_n, wave_gen_1_s0_translator:reset, wave_gen_1_s0_translator_avalon_universal_slave_0_agent:reset, wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, wave_gen_2:reset_n, wave_gen_2_s0_translator:reset, wave_gen_2_s0_translator_avalon_universal_slave_0_agent:reset, wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_002_reset_out_reset;                                                                 // rst_controller_002:reset_out -> ddr2:soft_reset_n
	wire          rst_controller_003_reset_out_reset;                                                                 // rst_controller_003:reset_out -> ddr2:global_reset_n
	wire          rst_controller_004_reset_out_reset;                                                                 // rst_controller_004:reset_out -> [altpll_0:reset, altpll_0_pll_slave_translator:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:out_reset, crosser_003:in_reset, id_router_006:reset, rsp_xbar_demux_006:reset]
	wire          rst_controller_005_reset_out_reset;                                                                 // rst_controller_005:reset_out -> [addr_router_005:reset, cmd_xbar_demux_005:reset, cpu_ddr2_clock_bridge:m0_reset, cpu_ddr2_clock_bridge_m0_translator:reset, cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                    // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                          // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                  // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire   [99:0] cmd_xbar_demux_src0_data;                                                                           // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire    [5:0] cmd_xbar_demux_src0_channel;                                                                        // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                          // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                    // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                          // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                  // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire   [99:0] cmd_xbar_demux_src1_data;                                                                           // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire    [5:0] cmd_xbar_demux_src1_channel;                                                                        // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                          // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                    // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                          // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                  // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire   [99:0] cmd_xbar_demux_src2_data;                                                                           // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire    [5:0] cmd_xbar_demux_src2_channel;                                                                        // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                          // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_src3_endofpacket;                                                                    // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                          // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                  // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire   [99:0] cmd_xbar_demux_src3_data;                                                                           // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire    [5:0] cmd_xbar_demux_src3_channel;                                                                        // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_src3_ready;                                                                          // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                      // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                              // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire   [99:0] cmd_xbar_demux_001_src0_data;                                                                       // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire    [5:0] cmd_xbar_demux_001_src0_channel;                                                                    // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                      // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                      // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                              // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire   [99:0] cmd_xbar_demux_001_src1_data;                                                                       // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire    [5:0] cmd_xbar_demux_001_src1_channel;                                                                    // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                      // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                      // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                              // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire   [99:0] cmd_xbar_demux_001_src2_data;                                                                       // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire    [5:0] cmd_xbar_demux_001_src2_channel;                                                                    // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                      // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                      // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                              // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire   [99:0] cmd_xbar_demux_001_src3_data;                                                                       // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire    [5:0] cmd_xbar_demux_001_src3_channel;                                                                    // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                      // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                // cmd_xbar_demux_001:src4_endofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                      // cmd_xbar_demux_001:src4_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                              // cmd_xbar_demux_001:src4_startofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [99:0] cmd_xbar_demux_001_src4_data;                                                                       // cmd_xbar_demux_001:src4_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_demux_001_src4_channel;                                                                    // cmd_xbar_demux_001:src4_channel -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                // cmd_xbar_demux_001:src5_endofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                      // cmd_xbar_demux_001:src5_valid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                              // cmd_xbar_demux_001:src5_startofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [99:0] cmd_xbar_demux_001_src5_data;                                                                       // cmd_xbar_demux_001:src5_data -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_demux_001_src5_channel;                                                                    // cmd_xbar_demux_001:src5_channel -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_003:sink2_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                      // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_003:sink2_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                              // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_003:sink2_startofpacket
	wire   [99:0] cmd_xbar_demux_002_src0_data;                                                                       // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_003:sink2_data
	wire    [5:0] cmd_xbar_demux_002_src0_channel;                                                                    // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_003:sink2_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                      // cmd_xbar_mux_003:sink2_ready -> cmd_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                    // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                          // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                  // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire   [99:0] rsp_xbar_demux_src0_data;                                                                           // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [5:0] rsp_xbar_demux_src0_channel;                                                                        // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                          // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                    // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                          // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                  // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire   [99:0] rsp_xbar_demux_src1_data;                                                                           // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire    [5:0] rsp_xbar_demux_src1_channel;                                                                        // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                          // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                      // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                              // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire   [99:0] rsp_xbar_demux_001_src0_data;                                                                       // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [5:0] rsp_xbar_demux_001_src0_channel;                                                                    // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                      // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                      // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                              // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire   [99:0] rsp_xbar_demux_001_src1_data;                                                                       // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire    [5:0] rsp_xbar_demux_001_src1_channel;                                                                    // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                      // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                      // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                              // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire   [99:0] rsp_xbar_demux_002_src0_data;                                                                       // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire    [5:0] rsp_xbar_demux_002_src0_channel;                                                                    // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                      // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                      // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                              // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire   [99:0] rsp_xbar_demux_002_src1_data;                                                                       // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire    [5:0] rsp_xbar_demux_002_src1_channel;                                                                    // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                      // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                      // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                              // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire   [99:0] rsp_xbar_demux_003_src0_data;                                                                       // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire    [5:0] rsp_xbar_demux_003_src0_channel;                                                                    // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                      // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                                // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                      // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                              // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire   [99:0] rsp_xbar_demux_003_src1_data;                                                                       // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire    [5:0] rsp_xbar_demux_003_src1_channel;                                                                    // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                      // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_003_src2_endofpacket;                                                                // rsp_xbar_demux_003:src2_endofpacket -> dma_0_read_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_003_src2_valid;                                                                      // rsp_xbar_demux_003:src2_valid -> dma_0_read_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_003_src2_startofpacket;                                                              // rsp_xbar_demux_003:src2_startofpacket -> dma_0_read_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [99:0] rsp_xbar_demux_003_src2_data;                                                                       // rsp_xbar_demux_003:src2_data -> dma_0_read_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] rsp_xbar_demux_003_src2_channel;                                                                    // rsp_xbar_demux_003:src2_channel -> dma_0_read_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                      // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                              // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire   [99:0] rsp_xbar_demux_004_src0_data;                                                                       // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire    [5:0] rsp_xbar_demux_004_src0_channel;                                                                    // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                      // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                      // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                              // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire   [99:0] rsp_xbar_demux_005_src0_data;                                                                       // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire    [5:0] rsp_xbar_demux_005_src0_channel;                                                                    // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                      // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                        // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                      // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire   [99:0] limiter_cmd_src_data;                                                                               // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire    [5:0] limiter_cmd_src_channel;                                                                            // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                              // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                       // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                             // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                     // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire   [99:0] rsp_xbar_mux_src_data;                                                                              // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire    [5:0] rsp_xbar_mux_src_channel;                                                                           // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                             // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                    // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                          // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                  // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire   [99:0] addr_router_001_src_data;                                                                           // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire    [5:0] addr_router_001_src_channel;                                                                        // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                          // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                   // rsp_xbar_mux_001:src_endofpacket -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                         // rsp_xbar_mux_001:src_valid -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                 // rsp_xbar_mux_001:src_startofpacket -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [99:0] rsp_xbar_mux_001_src_data;                                                                          // rsp_xbar_mux_001:src_data -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] rsp_xbar_mux_001_src_channel;                                                                       // rsp_xbar_mux_001:src_channel -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                         // nios2_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          addr_router_002_src_endofpacket;                                                                    // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                          // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                  // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire   [99:0] addr_router_002_src_data;                                                                           // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire    [5:0] addr_router_002_src_channel;                                                                        // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                          // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_demux_003_src2_ready;                                                                      // dma_0_read_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_003:src2_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                       // cmd_xbar_mux:src_endofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                             // cmd_xbar_mux:src_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                     // cmd_xbar_mux:src_startofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [99:0] cmd_xbar_mux_src_data;                                                                              // cmd_xbar_mux:src_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_mux_src_channel;                                                                           // cmd_xbar_mux:src_channel -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                             // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                          // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                        // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire   [99:0] id_router_src_data;                                                                                 // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [5:0] id_router_src_channel;                                                                              // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                   // cmd_xbar_mux_001:src_endofpacket -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                         // cmd_xbar_mux_001:src_valid -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                 // cmd_xbar_mux_001:src_startofpacket -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [99:0] cmd_xbar_mux_001_src_data;                                                                          // cmd_xbar_mux_001:src_data -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_mux_001_src_channel;                                                                       // cmd_xbar_mux_001:src_channel -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                         // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                      // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                            // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                    // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire   [99:0] id_router_001_src_data;                                                                             // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [5:0] id_router_001_src_channel;                                                                          // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                            // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                   // cmd_xbar_mux_002:src_endofpacket -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                         // cmd_xbar_mux_002:src_valid -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                 // cmd_xbar_mux_002:src_startofpacket -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [99:0] cmd_xbar_mux_002_src_data;                                                                          // cmd_xbar_mux_002:src_data -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_mux_002_src_channel;                                                                       // cmd_xbar_mux_002:src_channel -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                         // onchip_ram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                      // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                            // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                    // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire   [99:0] id_router_002_src_data;                                                                             // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [5:0] id_router_002_src_channel;                                                                          // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                            // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                   // cmd_xbar_mux_003:src_endofpacket -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                         // cmd_xbar_mux_003:src_valid -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                 // cmd_xbar_mux_003:src_startofpacket -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [99:0] cmd_xbar_mux_003_src_data;                                                                          // cmd_xbar_mux_003:src_data -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_mux_003_src_channel;                                                                       // cmd_xbar_mux_003:src_channel -> cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                         // cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire          id_router_003_src_endofpacket;                                                                      // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                            // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                    // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire   [99:0] id_router_003_src_data;                                                                             // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [5:0] id_router_003_src_channel;                                                                          // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                            // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                      // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_004_src_endofpacket;                                                                      // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                            // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                    // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire   [99:0] id_router_004_src_data;                                                                             // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire    [5:0] id_router_004_src_channel;                                                                          // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                            // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_001_src5_ready;                                                                      // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire          id_router_005_src_endofpacket;                                                                      // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                            // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                    // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire   [99:0] id_router_005_src_data;                                                                             // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire    [5:0] id_router_005_src_channel;                                                                          // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                            // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_003_src1_endofpacket;                                                                // cmd_xbar_demux_003:src1_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src1_valid;                                                                      // cmd_xbar_demux_003:src1_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src1_startofpacket;                                                              // cmd_xbar_demux_003:src1_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src1_data;                                                                       // cmd_xbar_demux_003:src1_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src1_channel;                                                                    // cmd_xbar_demux_003:src1_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src2_endofpacket;                                                                // cmd_xbar_demux_003:src2_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src2_valid;                                                                      // cmd_xbar_demux_003:src2_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src2_startofpacket;                                                              // cmd_xbar_demux_003:src2_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src2_data;                                                                       // cmd_xbar_demux_003:src2_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src2_channel;                                                                    // cmd_xbar_demux_003:src2_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src3_endofpacket;                                                                // cmd_xbar_demux_003:src3_endofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src3_valid;                                                                      // cmd_xbar_demux_003:src3_valid -> systimer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src3_startofpacket;                                                              // cmd_xbar_demux_003:src3_startofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src3_data;                                                                       // cmd_xbar_demux_003:src3_data -> systimer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src3_channel;                                                                    // cmd_xbar_demux_003:src3_channel -> systimer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src4_endofpacket;                                                                // cmd_xbar_demux_003:src4_endofpacket -> pio_key_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src4_valid;                                                                      // cmd_xbar_demux_003:src4_valid -> pio_key_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src4_startofpacket;                                                              // cmd_xbar_demux_003:src4_startofpacket -> pio_key_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src4_data;                                                                       // cmd_xbar_demux_003:src4_data -> pio_key_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src4_channel;                                                                    // cmd_xbar_demux_003:src4_channel -> pio_key_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src5_endofpacket;                                                                // cmd_xbar_demux_003:src5_endofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src5_valid;                                                                      // cmd_xbar_demux_003:src5_valid -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src5_startofpacket;                                                              // cmd_xbar_demux_003:src5_startofpacket -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src5_data;                                                                       // cmd_xbar_demux_003:src5_data -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src5_channel;                                                                    // cmd_xbar_demux_003:src5_channel -> spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src6_endofpacket;                                                                // cmd_xbar_demux_003:src6_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src6_valid;                                                                      // cmd_xbar_demux_003:src6_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src6_startofpacket;                                                              // cmd_xbar_demux_003:src6_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src6_data;                                                                       // cmd_xbar_demux_003:src6_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src6_channel;                                                                    // cmd_xbar_demux_003:src6_channel -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src7_endofpacket;                                                                // cmd_xbar_demux_003:src7_endofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src7_valid;                                                                      // cmd_xbar_demux_003:src7_valid -> pio_led_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src7_startofpacket;                                                              // cmd_xbar_demux_003:src7_startofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src7_data;                                                                       // cmd_xbar_demux_003:src7_data -> pio_led_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src7_channel;                                                                    // cmd_xbar_demux_003:src7_channel -> pio_led_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src8_endofpacket;                                                                // cmd_xbar_demux_003:src8_endofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src8_valid;                                                                      // cmd_xbar_demux_003:src8_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src8_startofpacket;                                                              // cmd_xbar_demux_003:src8_startofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src8_data;                                                                       // cmd_xbar_demux_003:src8_data -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src8_channel;                                                                    // cmd_xbar_demux_003:src8_channel -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src9_endofpacket;                                                                // cmd_xbar_demux_003:src9_endofpacket -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src9_valid;                                                                      // cmd_xbar_demux_003:src9_valid -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src9_startofpacket;                                                              // cmd_xbar_demux_003:src9_startofpacket -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src9_data;                                                                       // cmd_xbar_demux_003:src9_data -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src9_channel;                                                                    // cmd_xbar_demux_003:src9_channel -> spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src10_endofpacket;                                                               // cmd_xbar_demux_003:src10_endofpacket -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src10_valid;                                                                     // cmd_xbar_demux_003:src10_valid -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src10_startofpacket;                                                             // cmd_xbar_demux_003:src10_startofpacket -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src10_data;                                                                      // cmd_xbar_demux_003:src10_data -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src10_channel;                                                                   // cmd_xbar_demux_003:src10_channel -> ad9245_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src11_endofpacket;                                                               // cmd_xbar_demux_003:src11_endofpacket -> clk_gen_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src11_valid;                                                                     // cmd_xbar_demux_003:src11_valid -> clk_gen_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src11_startofpacket;                                                             // cmd_xbar_demux_003:src11_startofpacket -> clk_gen_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src11_data;                                                                      // cmd_xbar_demux_003:src11_data -> clk_gen_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src11_channel;                                                                   // cmd_xbar_demux_003:src11_channel -> clk_gen_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src12_endofpacket;                                                               // cmd_xbar_demux_003:src12_endofpacket -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src12_valid;                                                                     // cmd_xbar_demux_003:src12_valid -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src12_startofpacket;                                                             // cmd_xbar_demux_003:src12_startofpacket -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src12_data;                                                                      // cmd_xbar_demux_003:src12_data -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src12_channel;                                                                   // cmd_xbar_demux_003:src12_channel -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src13_endofpacket;                                                               // cmd_xbar_demux_003:src13_endofpacket -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src13_valid;                                                                     // cmd_xbar_demux_003:src13_valid -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src13_startofpacket;                                                             // cmd_xbar_demux_003:src13_startofpacket -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src13_data;                                                                      // cmd_xbar_demux_003:src13_data -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src13_channel;                                                                   // cmd_xbar_demux_003:src13_channel -> spi_master_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src14_endofpacket;                                                               // cmd_xbar_demux_003:src14_endofpacket -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src14_valid;                                                                     // cmd_xbar_demux_003:src14_valid -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src14_startofpacket;                                                             // cmd_xbar_demux_003:src14_startofpacket -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src14_data;                                                                      // cmd_xbar_demux_003:src14_data -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src14_channel;                                                                   // cmd_xbar_demux_003:src14_channel -> ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src15_endofpacket;                                                               // cmd_xbar_demux_003:src15_endofpacket -> cmd_xbar_mux_021:sink0_endofpacket
	wire          cmd_xbar_demux_003_src15_valid;                                                                     // cmd_xbar_demux_003:src15_valid -> cmd_xbar_mux_021:sink0_valid
	wire          cmd_xbar_demux_003_src15_startofpacket;                                                             // cmd_xbar_demux_003:src15_startofpacket -> cmd_xbar_mux_021:sink0_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src15_data;                                                                      // cmd_xbar_demux_003:src15_data -> cmd_xbar_mux_021:sink0_data
	wire   [23:0] cmd_xbar_demux_003_src15_channel;                                                                   // cmd_xbar_demux_003:src15_channel -> cmd_xbar_mux_021:sink0_channel
	wire          cmd_xbar_demux_003_src15_ready;                                                                     // cmd_xbar_mux_021:sink0_ready -> cmd_xbar_demux_003:src15_ready
	wire          cmd_xbar_demux_003_src16_endofpacket;                                                               // cmd_xbar_demux_003:src16_endofpacket -> cmd_xbar_mux_022:sink0_endofpacket
	wire          cmd_xbar_demux_003_src16_valid;                                                                     // cmd_xbar_demux_003:src16_valid -> cmd_xbar_mux_022:sink0_valid
	wire          cmd_xbar_demux_003_src16_startofpacket;                                                             // cmd_xbar_demux_003:src16_startofpacket -> cmd_xbar_mux_022:sink0_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src16_data;                                                                      // cmd_xbar_demux_003:src16_data -> cmd_xbar_mux_022:sink0_data
	wire   [23:0] cmd_xbar_demux_003_src16_channel;                                                                   // cmd_xbar_demux_003:src16_channel -> cmd_xbar_mux_022:sink0_channel
	wire          cmd_xbar_demux_003_src16_ready;                                                                     // cmd_xbar_mux_022:sink0_ready -> cmd_xbar_demux_003:src16_ready
	wire          cmd_xbar_demux_003_src17_endofpacket;                                                               // cmd_xbar_demux_003:src17_endofpacket -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src17_valid;                                                                     // cmd_xbar_demux_003:src17_valid -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src17_startofpacket;                                                             // cmd_xbar_demux_003:src17_startofpacket -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src17_data;                                                                      // cmd_xbar_demux_003:src17_data -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src17_channel;                                                                   // cmd_xbar_demux_003:src17_channel -> dac2904_2_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src18_endofpacket;                                                               // cmd_xbar_demux_003:src18_endofpacket -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src18_valid;                                                                     // cmd_xbar_demux_003:src18_valid -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src18_startofpacket;                                                             // cmd_xbar_demux_003:src18_startofpacket -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src18_data;                                                                      // cmd_xbar_demux_003:src18_data -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src18_channel;                                                                   // cmd_xbar_demux_003:src18_channel -> dac2904_3_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src19_endofpacket;                                                               // cmd_xbar_demux_003:src19_endofpacket -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src19_valid;                                                                     // cmd_xbar_demux_003:src19_valid -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src19_startofpacket;                                                             // cmd_xbar_demux_003:src19_startofpacket -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src19_data;                                                                      // cmd_xbar_demux_003:src19_data -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src19_channel;                                                                   // cmd_xbar_demux_003:src19_channel -> dac2904_4_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src20_endofpacket;                                                               // cmd_xbar_demux_003:src20_endofpacket -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src20_valid;                                                                     // cmd_xbar_demux_003:src20_valid -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src20_startofpacket;                                                             // cmd_xbar_demux_003:src20_startofpacket -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src20_data;                                                                      // cmd_xbar_demux_003:src20_data -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src20_channel;                                                                   // cmd_xbar_demux_003:src20_channel -> wave_gen_0_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src21_endofpacket;                                                               // cmd_xbar_demux_003:src21_endofpacket -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src21_valid;                                                                     // cmd_xbar_demux_003:src21_valid -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src21_startofpacket;                                                             // cmd_xbar_demux_003:src21_startofpacket -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src21_data;                                                                      // cmd_xbar_demux_003:src21_data -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src21_channel;                                                                   // cmd_xbar_demux_003:src21_channel -> demodulation_0_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src22_endofpacket;                                                               // cmd_xbar_demux_003:src22_endofpacket -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src22_valid;                                                                     // cmd_xbar_demux_003:src22_valid -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src22_startofpacket;                                                             // cmd_xbar_demux_003:src22_startofpacket -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src22_data;                                                                      // cmd_xbar_demux_003:src22_data -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src22_channel;                                                                   // cmd_xbar_demux_003:src22_channel -> wave_gen_1_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src23_endofpacket;                                                               // cmd_xbar_demux_003:src23_endofpacket -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src23_valid;                                                                     // cmd_xbar_demux_003:src23_valid -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src23_startofpacket;                                                             // cmd_xbar_demux_003:src23_startofpacket -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src23_data;                                                                      // cmd_xbar_demux_003:src23_data -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_demux_003_src23_channel;                                                                   // cmd_xbar_demux_003:src23_channel -> wave_gen_2_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_003:sink1_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                      // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_003:sink1_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                              // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_003:sink1_startofpacket
	wire   [84:0] rsp_xbar_demux_007_src0_data;                                                                       // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_003:sink1_data
	wire   [23:0] rsp_xbar_demux_007_src0_channel;                                                                    // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_003:sink1_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                      // rsp_xbar_mux_003:sink1_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_003:sink2_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                      // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_003:sink2_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                              // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_003:sink2_startofpacket
	wire   [84:0] rsp_xbar_demux_008_src0_data;                                                                       // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_003:sink2_data
	wire   [23:0] rsp_xbar_demux_008_src0_channel;                                                                    // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_003:sink2_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                      // rsp_xbar_mux_003:sink2_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_003:sink3_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                      // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_003:sink3_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                              // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_003:sink3_startofpacket
	wire   [84:0] rsp_xbar_demux_009_src0_data;                                                                       // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_003:sink3_data
	wire   [23:0] rsp_xbar_demux_009_src0_channel;                                                                    // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_003:sink3_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                      // rsp_xbar_mux_003:sink3_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_003:sink4_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                      // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_003:sink4_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                              // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_003:sink4_startofpacket
	wire   [84:0] rsp_xbar_demux_010_src0_data;                                                                       // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_003:sink4_data
	wire   [23:0] rsp_xbar_demux_010_src0_channel;                                                                    // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_003:sink4_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                      // rsp_xbar_mux_003:sink4_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_003:sink5_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                      // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_003:sink5_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                              // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_003:sink5_startofpacket
	wire   [84:0] rsp_xbar_demux_011_src0_data;                                                                       // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_003:sink5_data
	wire   [23:0] rsp_xbar_demux_011_src0_channel;                                                                    // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_003:sink5_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                      // rsp_xbar_mux_003:sink5_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_003:sink6_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                      // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_003:sink6_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                              // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_003:sink6_startofpacket
	wire   [84:0] rsp_xbar_demux_012_src0_data;                                                                       // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_003:sink6_data
	wire   [23:0] rsp_xbar_demux_012_src0_channel;                                                                    // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_003:sink6_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                      // rsp_xbar_mux_003:sink6_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_003:sink7_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                      // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_003:sink7_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                              // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_003:sink7_startofpacket
	wire   [84:0] rsp_xbar_demux_013_src0_data;                                                                       // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_003:sink7_data
	wire   [23:0] rsp_xbar_demux_013_src0_channel;                                                                    // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_003:sink7_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                      // rsp_xbar_mux_003:sink7_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_003:sink8_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                      // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_003:sink8_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                              // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_003:sink8_startofpacket
	wire   [84:0] rsp_xbar_demux_014_src0_data;                                                                       // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_003:sink8_data
	wire   [23:0] rsp_xbar_demux_014_src0_channel;                                                                    // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_003:sink8_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                      // rsp_xbar_mux_003:sink8_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_003:sink9_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                      // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_003:sink9_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                              // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_003:sink9_startofpacket
	wire   [84:0] rsp_xbar_demux_015_src0_data;                                                                       // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_003:sink9_data
	wire   [23:0] rsp_xbar_demux_015_src0_channel;                                                                    // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_003:sink9_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                      // rsp_xbar_mux_003:sink9_ready -> rsp_xbar_demux_015:src0_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                                // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_003:sink10_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                      // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_003:sink10_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                              // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_003:sink10_startofpacket
	wire   [84:0] rsp_xbar_demux_016_src0_data;                                                                       // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_003:sink10_data
	wire   [23:0] rsp_xbar_demux_016_src0_channel;                                                                    // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_003:sink10_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                      // rsp_xbar_mux_003:sink10_ready -> rsp_xbar_demux_016:src0_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                                // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_003:sink11_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                      // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_003:sink11_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                              // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_003:sink11_startofpacket
	wire   [84:0] rsp_xbar_demux_017_src0_data;                                                                       // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_003:sink11_data
	wire   [23:0] rsp_xbar_demux_017_src0_channel;                                                                    // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_003:sink11_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                      // rsp_xbar_mux_003:sink11_ready -> rsp_xbar_demux_017:src0_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                                // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_003:sink12_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                      // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_003:sink12_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                              // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_003:sink12_startofpacket
	wire   [84:0] rsp_xbar_demux_018_src0_data;                                                                       // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_003:sink12_data
	wire   [23:0] rsp_xbar_demux_018_src0_channel;                                                                    // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_003:sink12_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                      // rsp_xbar_mux_003:sink12_ready -> rsp_xbar_demux_018:src0_ready
	wire          rsp_xbar_demux_019_src0_endofpacket;                                                                // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_003:sink13_endofpacket
	wire          rsp_xbar_demux_019_src0_valid;                                                                      // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_003:sink13_valid
	wire          rsp_xbar_demux_019_src0_startofpacket;                                                              // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_003:sink13_startofpacket
	wire   [84:0] rsp_xbar_demux_019_src0_data;                                                                       // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_003:sink13_data
	wire   [23:0] rsp_xbar_demux_019_src0_channel;                                                                    // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_003:sink13_channel
	wire          rsp_xbar_demux_019_src0_ready;                                                                      // rsp_xbar_mux_003:sink13_ready -> rsp_xbar_demux_019:src0_ready
	wire          rsp_xbar_demux_020_src0_endofpacket;                                                                // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_003:sink14_endofpacket
	wire          rsp_xbar_demux_020_src0_valid;                                                                      // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_003:sink14_valid
	wire          rsp_xbar_demux_020_src0_startofpacket;                                                              // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_003:sink14_startofpacket
	wire   [84:0] rsp_xbar_demux_020_src0_data;                                                                       // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_003:sink14_data
	wire   [23:0] rsp_xbar_demux_020_src0_channel;                                                                    // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_003:sink14_channel
	wire          rsp_xbar_demux_020_src0_ready;                                                                      // rsp_xbar_mux_003:sink14_ready -> rsp_xbar_demux_020:src0_ready
	wire          rsp_xbar_demux_021_src0_endofpacket;                                                                // rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_003:sink15_endofpacket
	wire          rsp_xbar_demux_021_src0_valid;                                                                      // rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_003:sink15_valid
	wire          rsp_xbar_demux_021_src0_startofpacket;                                                              // rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_003:sink15_startofpacket
	wire   [84:0] rsp_xbar_demux_021_src0_data;                                                                       // rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_003:sink15_data
	wire   [23:0] rsp_xbar_demux_021_src0_channel;                                                                    // rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_003:sink15_channel
	wire          rsp_xbar_demux_021_src0_ready;                                                                      // rsp_xbar_mux_003:sink15_ready -> rsp_xbar_demux_021:src0_ready
	wire          rsp_xbar_demux_022_src0_endofpacket;                                                                // rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux_003:sink16_endofpacket
	wire          rsp_xbar_demux_022_src0_valid;                                                                      // rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux_003:sink16_valid
	wire          rsp_xbar_demux_022_src0_startofpacket;                                                              // rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux_003:sink16_startofpacket
	wire   [84:0] rsp_xbar_demux_022_src0_data;                                                                       // rsp_xbar_demux_022:src0_data -> rsp_xbar_mux_003:sink16_data
	wire   [23:0] rsp_xbar_demux_022_src0_channel;                                                                    // rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux_003:sink16_channel
	wire          rsp_xbar_demux_022_src0_ready;                                                                      // rsp_xbar_mux_003:sink16_ready -> rsp_xbar_demux_022:src0_ready
	wire          rsp_xbar_demux_023_src0_endofpacket;                                                                // rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux_003:sink17_endofpacket
	wire          rsp_xbar_demux_023_src0_valid;                                                                      // rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux_003:sink17_valid
	wire          rsp_xbar_demux_023_src0_startofpacket;                                                              // rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux_003:sink17_startofpacket
	wire   [84:0] rsp_xbar_demux_023_src0_data;                                                                       // rsp_xbar_demux_023:src0_data -> rsp_xbar_mux_003:sink17_data
	wire   [23:0] rsp_xbar_demux_023_src0_channel;                                                                    // rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux_003:sink17_channel
	wire          rsp_xbar_demux_023_src0_ready;                                                                      // rsp_xbar_mux_003:sink17_ready -> rsp_xbar_demux_023:src0_ready
	wire          rsp_xbar_demux_024_src0_endofpacket;                                                                // rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux_003:sink18_endofpacket
	wire          rsp_xbar_demux_024_src0_valid;                                                                      // rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux_003:sink18_valid
	wire          rsp_xbar_demux_024_src0_startofpacket;                                                              // rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux_003:sink18_startofpacket
	wire   [84:0] rsp_xbar_demux_024_src0_data;                                                                       // rsp_xbar_demux_024:src0_data -> rsp_xbar_mux_003:sink18_data
	wire   [23:0] rsp_xbar_demux_024_src0_channel;                                                                    // rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux_003:sink18_channel
	wire          rsp_xbar_demux_024_src0_ready;                                                                      // rsp_xbar_mux_003:sink18_ready -> rsp_xbar_demux_024:src0_ready
	wire          rsp_xbar_demux_025_src0_endofpacket;                                                                // rsp_xbar_demux_025:src0_endofpacket -> rsp_xbar_mux_003:sink19_endofpacket
	wire          rsp_xbar_demux_025_src0_valid;                                                                      // rsp_xbar_demux_025:src0_valid -> rsp_xbar_mux_003:sink19_valid
	wire          rsp_xbar_demux_025_src0_startofpacket;                                                              // rsp_xbar_demux_025:src0_startofpacket -> rsp_xbar_mux_003:sink19_startofpacket
	wire   [84:0] rsp_xbar_demux_025_src0_data;                                                                       // rsp_xbar_demux_025:src0_data -> rsp_xbar_mux_003:sink19_data
	wire   [23:0] rsp_xbar_demux_025_src0_channel;                                                                    // rsp_xbar_demux_025:src0_channel -> rsp_xbar_mux_003:sink19_channel
	wire          rsp_xbar_demux_025_src0_ready;                                                                      // rsp_xbar_mux_003:sink19_ready -> rsp_xbar_demux_025:src0_ready
	wire          rsp_xbar_demux_026_src0_endofpacket;                                                                // rsp_xbar_demux_026:src0_endofpacket -> rsp_xbar_mux_003:sink20_endofpacket
	wire          rsp_xbar_demux_026_src0_valid;                                                                      // rsp_xbar_demux_026:src0_valid -> rsp_xbar_mux_003:sink20_valid
	wire          rsp_xbar_demux_026_src0_startofpacket;                                                              // rsp_xbar_demux_026:src0_startofpacket -> rsp_xbar_mux_003:sink20_startofpacket
	wire   [84:0] rsp_xbar_demux_026_src0_data;                                                                       // rsp_xbar_demux_026:src0_data -> rsp_xbar_mux_003:sink20_data
	wire   [23:0] rsp_xbar_demux_026_src0_channel;                                                                    // rsp_xbar_demux_026:src0_channel -> rsp_xbar_mux_003:sink20_channel
	wire          rsp_xbar_demux_026_src0_ready;                                                                      // rsp_xbar_mux_003:sink20_ready -> rsp_xbar_demux_026:src0_ready
	wire          rsp_xbar_demux_027_src0_endofpacket;                                                                // rsp_xbar_demux_027:src0_endofpacket -> rsp_xbar_mux_003:sink21_endofpacket
	wire          rsp_xbar_demux_027_src0_valid;                                                                      // rsp_xbar_demux_027:src0_valid -> rsp_xbar_mux_003:sink21_valid
	wire          rsp_xbar_demux_027_src0_startofpacket;                                                              // rsp_xbar_demux_027:src0_startofpacket -> rsp_xbar_mux_003:sink21_startofpacket
	wire   [84:0] rsp_xbar_demux_027_src0_data;                                                                       // rsp_xbar_demux_027:src0_data -> rsp_xbar_mux_003:sink21_data
	wire   [23:0] rsp_xbar_demux_027_src0_channel;                                                                    // rsp_xbar_demux_027:src0_channel -> rsp_xbar_mux_003:sink21_channel
	wire          rsp_xbar_demux_027_src0_ready;                                                                      // rsp_xbar_mux_003:sink21_ready -> rsp_xbar_demux_027:src0_ready
	wire          rsp_xbar_demux_028_src0_endofpacket;                                                                // rsp_xbar_demux_028:src0_endofpacket -> rsp_xbar_mux_003:sink22_endofpacket
	wire          rsp_xbar_demux_028_src0_valid;                                                                      // rsp_xbar_demux_028:src0_valid -> rsp_xbar_mux_003:sink22_valid
	wire          rsp_xbar_demux_028_src0_startofpacket;                                                              // rsp_xbar_demux_028:src0_startofpacket -> rsp_xbar_mux_003:sink22_startofpacket
	wire   [84:0] rsp_xbar_demux_028_src0_data;                                                                       // rsp_xbar_demux_028:src0_data -> rsp_xbar_mux_003:sink22_data
	wire   [23:0] rsp_xbar_demux_028_src0_channel;                                                                    // rsp_xbar_demux_028:src0_channel -> rsp_xbar_mux_003:sink22_channel
	wire          rsp_xbar_demux_028_src0_ready;                                                                      // rsp_xbar_mux_003:sink22_ready -> rsp_xbar_demux_028:src0_ready
	wire          rsp_xbar_demux_029_src0_endofpacket;                                                                // rsp_xbar_demux_029:src0_endofpacket -> rsp_xbar_mux_003:sink23_endofpacket
	wire          rsp_xbar_demux_029_src0_valid;                                                                      // rsp_xbar_demux_029:src0_valid -> rsp_xbar_mux_003:sink23_valid
	wire          rsp_xbar_demux_029_src0_startofpacket;                                                              // rsp_xbar_demux_029:src0_startofpacket -> rsp_xbar_mux_003:sink23_startofpacket
	wire   [84:0] rsp_xbar_demux_029_src0_data;                                                                       // rsp_xbar_demux_029:src0_data -> rsp_xbar_mux_003:sink23_data
	wire   [23:0] rsp_xbar_demux_029_src0_channel;                                                                    // rsp_xbar_demux_029:src0_channel -> rsp_xbar_mux_003:sink23_channel
	wire          rsp_xbar_demux_029_src0_ready;                                                                      // rsp_xbar_mux_003:sink23_ready -> rsp_xbar_demux_029:src0_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                    // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                  // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire   [84:0] limiter_001_cmd_src_data;                                                                           // limiter_001:cmd_src_data -> cmd_xbar_demux_003:sink_data
	wire   [23:0] limiter_001_cmd_src_channel;                                                                        // limiter_001:cmd_src_channel -> cmd_xbar_demux_003:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                          // cmd_xbar_demux_003:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_003_src_endofpacket;                                                                   // rsp_xbar_mux_003:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_003_src_valid;                                                                         // rsp_xbar_mux_003:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_003_src_startofpacket;                                                                 // rsp_xbar_mux_003:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire   [84:0] rsp_xbar_mux_003_src_data;                                                                          // rsp_xbar_mux_003:src_data -> limiter_001:rsp_sink_data
	wire   [23:0] rsp_xbar_mux_003_src_channel;                                                                       // rsp_xbar_mux_003:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_003_src_ready;                                                                         // limiter_001:rsp_sink_ready -> rsp_xbar_mux_003:src_ready
	wire          addr_router_004_src_endofpacket;                                                                    // addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          addr_router_004_src_valid;                                                                          // addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	wire          addr_router_004_src_startofpacket;                                                                  // addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire   [84:0] addr_router_004_src_data;                                                                           // addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	wire   [23:0] addr_router_004_src_channel;                                                                        // addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	wire          addr_router_004_src_ready;                                                                          // cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	wire          rsp_xbar_mux_004_src_endofpacket;                                                                   // rsp_xbar_mux_004:src_endofpacket -> dma_0_write_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_004_src_valid;                                                                         // rsp_xbar_mux_004:src_valid -> dma_0_write_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_004_src_startofpacket;                                                                 // rsp_xbar_mux_004:src_startofpacket -> dma_0_write_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [84:0] rsp_xbar_mux_004_src_data;                                                                          // rsp_xbar_mux_004:src_data -> dma_0_write_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [23:0] rsp_xbar_mux_004_src_channel;                                                                       // rsp_xbar_mux_004:src_channel -> dma_0_write_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_004_src_ready;                                                                         // dma_0_write_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_004:src_ready
	wire          crosser_out_ready;                                                                                  // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire          id_router_006_src_endofpacket;                                                                      // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                            // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                    // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire   [84:0] id_router_006_src_data;                                                                             // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [23:0] id_router_006_src_channel;                                                                          // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                            // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_003_src1_ready;                                                                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src1_ready
	wire          id_router_007_src_endofpacket;                                                                      // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                            // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                    // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire   [84:0] id_router_007_src_data;                                                                             // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [23:0] id_router_007_src_channel;                                                                          // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                            // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_003_src2_ready;                                                                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src2_ready
	wire          id_router_008_src_endofpacket;                                                                      // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                            // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                    // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire   [84:0] id_router_008_src_data;                                                                             // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [23:0] id_router_008_src_channel;                                                                          // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                            // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_003_src3_ready;                                                                      // systimer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src3_ready
	wire          id_router_009_src_endofpacket;                                                                      // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                            // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                    // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire   [84:0] id_router_009_src_data;                                                                             // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [23:0] id_router_009_src_channel;                                                                          // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                            // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_003_src4_ready;                                                                      // pio_key_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src4_ready
	wire          id_router_010_src_endofpacket;                                                                      // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                            // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                    // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire   [84:0] id_router_010_src_data;                                                                             // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [23:0] id_router_010_src_channel;                                                                          // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                            // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_003_src5_ready;                                                                      // spi_0_spi_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src5_ready
	wire          id_router_011_src_endofpacket;                                                                      // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                            // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                    // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire   [84:0] id_router_011_src_data;                                                                             // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [23:0] id_router_011_src_channel;                                                                          // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                            // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_003_src6_ready;                                                                      // uart_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src6_ready
	wire          id_router_012_src_endofpacket;                                                                      // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                            // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                    // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire   [84:0] id_router_012_src_data;                                                                             // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [23:0] id_router_012_src_channel;                                                                          // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                            // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_demux_003_src7_ready;                                                                      // pio_led_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src7_ready
	wire          id_router_013_src_endofpacket;                                                                      // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                            // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                    // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire   [84:0] id_router_013_src_data;                                                                             // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [23:0] id_router_013_src_channel;                                                                          // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                            // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_003_src8_ready;                                                                      // timestamp_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src8_ready
	wire          id_router_014_src_endofpacket;                                                                      // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                            // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                    // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire   [84:0] id_router_014_src_data;                                                                             // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [23:0] id_router_014_src_channel;                                                                          // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                            // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_003_src9_ready;                                                                      // spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src9_ready
	wire          id_router_015_src_endofpacket;                                                                      // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                            // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                    // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire   [84:0] id_router_015_src_data;                                                                             // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [23:0] id_router_015_src_channel;                                                                          // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                            // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_003_src10_ready;                                                                     // ad9245_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src10_ready
	wire          id_router_016_src_endofpacket;                                                                      // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                            // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                    // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire   [84:0] id_router_016_src_data;                                                                             // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [23:0] id_router_016_src_channel;                                                                          // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                            // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          cmd_xbar_demux_003_src11_ready;                                                                     // clk_gen_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src11_ready
	wire          id_router_017_src_endofpacket;                                                                      // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                            // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                    // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire   [84:0] id_router_017_src_data;                                                                             // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [23:0] id_router_017_src_channel;                                                                          // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                            // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          cmd_xbar_demux_003_src12_ready;                                                                     // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src12_ready
	wire          id_router_018_src_endofpacket;                                                                      // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                            // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                    // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire   [84:0] id_router_018_src_data;                                                                             // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire   [23:0] id_router_018_src_channel;                                                                          // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                            // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          cmd_xbar_demux_003_src13_ready;                                                                     // spi_master_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src13_ready
	wire          id_router_019_src_endofpacket;                                                                      // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire          id_router_019_src_valid;                                                                            // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire          id_router_019_src_startofpacket;                                                                    // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire   [84:0] id_router_019_src_data;                                                                             // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire   [23:0] id_router_019_src_channel;                                                                          // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire          id_router_019_src_ready;                                                                            // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire          cmd_xbar_demux_003_src14_ready;                                                                     // ad9266_spi_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src14_ready
	wire          id_router_020_src_endofpacket;                                                                      // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire          id_router_020_src_valid;                                                                            // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire          id_router_020_src_startofpacket;                                                                    // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire   [84:0] id_router_020_src_data;                                                                             // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire   [23:0] id_router_020_src_channel;                                                                          // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire          id_router_020_src_ready;                                                                            // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire          cmd_xbar_mux_021_src_endofpacket;                                                                   // cmd_xbar_mux_021:src_endofpacket -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_021_src_valid;                                                                         // cmd_xbar_mux_021:src_valid -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_021_src_startofpacket;                                                                 // cmd_xbar_mux_021:src_startofpacket -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_mux_021_src_data;                                                                          // cmd_xbar_mux_021:src_data -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_mux_021_src_channel;                                                                       // cmd_xbar_mux_021:src_channel -> ad9245_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_021_src_ready;                                                                         // ad9245_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_021:src_ready
	wire          id_router_021_src_endofpacket;                                                                      // id_router_021:src_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire          id_router_021_src_valid;                                                                            // id_router_021:src_valid -> rsp_xbar_demux_021:sink_valid
	wire          id_router_021_src_startofpacket;                                                                    // id_router_021:src_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire   [84:0] id_router_021_src_data;                                                                             // id_router_021:src_data -> rsp_xbar_demux_021:sink_data
	wire   [23:0] id_router_021_src_channel;                                                                          // id_router_021:src_channel -> rsp_xbar_demux_021:sink_channel
	wire          id_router_021_src_ready;                                                                            // rsp_xbar_demux_021:sink_ready -> id_router_021:src_ready
	wire          cmd_xbar_mux_022_src_endofpacket;                                                                   // cmd_xbar_mux_022:src_endofpacket -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_022_src_valid;                                                                         // cmd_xbar_mux_022:src_valid -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_022_src_startofpacket;                                                                 // cmd_xbar_mux_022:src_startofpacket -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] cmd_xbar_mux_022_src_data;                                                                          // cmd_xbar_mux_022:src_data -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] cmd_xbar_mux_022_src_channel;                                                                       // cmd_xbar_mux_022:src_channel -> dac2904_1_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_022_src_ready;                                                                         // dac2904_1_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_022:src_ready
	wire          id_router_022_src_endofpacket;                                                                      // id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire          id_router_022_src_valid;                                                                            // id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	wire          id_router_022_src_startofpacket;                                                                    // id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire   [84:0] id_router_022_src_data;                                                                             // id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	wire   [23:0] id_router_022_src_channel;                                                                          // id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	wire          id_router_022_src_ready;                                                                            // rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	wire          cmd_xbar_demux_003_src17_ready;                                                                     // dac2904_2_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src17_ready
	wire          id_router_023_src_endofpacket;                                                                      // id_router_023:src_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	wire          id_router_023_src_valid;                                                                            // id_router_023:src_valid -> rsp_xbar_demux_023:sink_valid
	wire          id_router_023_src_startofpacket;                                                                    // id_router_023:src_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	wire   [84:0] id_router_023_src_data;                                                                             // id_router_023:src_data -> rsp_xbar_demux_023:sink_data
	wire   [23:0] id_router_023_src_channel;                                                                          // id_router_023:src_channel -> rsp_xbar_demux_023:sink_channel
	wire          id_router_023_src_ready;                                                                            // rsp_xbar_demux_023:sink_ready -> id_router_023:src_ready
	wire          cmd_xbar_demux_003_src18_ready;                                                                     // dac2904_3_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src18_ready
	wire          id_router_024_src_endofpacket;                                                                      // id_router_024:src_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	wire          id_router_024_src_valid;                                                                            // id_router_024:src_valid -> rsp_xbar_demux_024:sink_valid
	wire          id_router_024_src_startofpacket;                                                                    // id_router_024:src_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	wire   [84:0] id_router_024_src_data;                                                                             // id_router_024:src_data -> rsp_xbar_demux_024:sink_data
	wire   [23:0] id_router_024_src_channel;                                                                          // id_router_024:src_channel -> rsp_xbar_demux_024:sink_channel
	wire          id_router_024_src_ready;                                                                            // rsp_xbar_demux_024:sink_ready -> id_router_024:src_ready
	wire          cmd_xbar_demux_003_src19_ready;                                                                     // dac2904_4_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src19_ready
	wire          id_router_025_src_endofpacket;                                                                      // id_router_025:src_endofpacket -> rsp_xbar_demux_025:sink_endofpacket
	wire          id_router_025_src_valid;                                                                            // id_router_025:src_valid -> rsp_xbar_demux_025:sink_valid
	wire          id_router_025_src_startofpacket;                                                                    // id_router_025:src_startofpacket -> rsp_xbar_demux_025:sink_startofpacket
	wire   [84:0] id_router_025_src_data;                                                                             // id_router_025:src_data -> rsp_xbar_demux_025:sink_data
	wire   [23:0] id_router_025_src_channel;                                                                          // id_router_025:src_channel -> rsp_xbar_demux_025:sink_channel
	wire          id_router_025_src_ready;                                                                            // rsp_xbar_demux_025:sink_ready -> id_router_025:src_ready
	wire          cmd_xbar_demux_003_src20_ready;                                                                     // wave_gen_0_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src20_ready
	wire          id_router_026_src_endofpacket;                                                                      // id_router_026:src_endofpacket -> rsp_xbar_demux_026:sink_endofpacket
	wire          id_router_026_src_valid;                                                                            // id_router_026:src_valid -> rsp_xbar_demux_026:sink_valid
	wire          id_router_026_src_startofpacket;                                                                    // id_router_026:src_startofpacket -> rsp_xbar_demux_026:sink_startofpacket
	wire   [84:0] id_router_026_src_data;                                                                             // id_router_026:src_data -> rsp_xbar_demux_026:sink_data
	wire   [23:0] id_router_026_src_channel;                                                                          // id_router_026:src_channel -> rsp_xbar_demux_026:sink_channel
	wire          id_router_026_src_ready;                                                                            // rsp_xbar_demux_026:sink_ready -> id_router_026:src_ready
	wire          cmd_xbar_demux_003_src21_ready;                                                                     // demodulation_0_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src21_ready
	wire          id_router_027_src_endofpacket;                                                                      // id_router_027:src_endofpacket -> rsp_xbar_demux_027:sink_endofpacket
	wire          id_router_027_src_valid;                                                                            // id_router_027:src_valid -> rsp_xbar_demux_027:sink_valid
	wire          id_router_027_src_startofpacket;                                                                    // id_router_027:src_startofpacket -> rsp_xbar_demux_027:sink_startofpacket
	wire   [84:0] id_router_027_src_data;                                                                             // id_router_027:src_data -> rsp_xbar_demux_027:sink_data
	wire   [23:0] id_router_027_src_channel;                                                                          // id_router_027:src_channel -> rsp_xbar_demux_027:sink_channel
	wire          id_router_027_src_ready;                                                                            // rsp_xbar_demux_027:sink_ready -> id_router_027:src_ready
	wire          cmd_xbar_demux_003_src22_ready;                                                                     // wave_gen_1_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src22_ready
	wire          id_router_028_src_endofpacket;                                                                      // id_router_028:src_endofpacket -> rsp_xbar_demux_028:sink_endofpacket
	wire          id_router_028_src_valid;                                                                            // id_router_028:src_valid -> rsp_xbar_demux_028:sink_valid
	wire          id_router_028_src_startofpacket;                                                                    // id_router_028:src_startofpacket -> rsp_xbar_demux_028:sink_startofpacket
	wire   [84:0] id_router_028_src_data;                                                                             // id_router_028:src_data -> rsp_xbar_demux_028:sink_data
	wire   [23:0] id_router_028_src_channel;                                                                          // id_router_028:src_channel -> rsp_xbar_demux_028:sink_channel
	wire          id_router_028_src_ready;                                                                            // rsp_xbar_demux_028:sink_ready -> id_router_028:src_ready
	wire          cmd_xbar_demux_003_src23_ready;                                                                     // wave_gen_2_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src23_ready
	wire          id_router_029_src_endofpacket;                                                                      // id_router_029:src_endofpacket -> rsp_xbar_demux_029:sink_endofpacket
	wire          id_router_029_src_valid;                                                                            // id_router_029:src_valid -> rsp_xbar_demux_029:sink_valid
	wire          id_router_029_src_startofpacket;                                                                    // id_router_029:src_startofpacket -> rsp_xbar_demux_029:sink_startofpacket
	wire   [84:0] id_router_029_src_data;                                                                             // id_router_029:src_data -> rsp_xbar_demux_029:sink_data
	wire   [23:0] id_router_029_src_channel;                                                                          // id_router_029:src_channel -> rsp_xbar_demux_029:sink_channel
	wire          id_router_029_src_ready;                                                                            // rsp_xbar_demux_029:sink_ready -> id_router_029:src_ready
	wire          cmd_xbar_demux_005_src0_endofpacket;                                                                // cmd_xbar_demux_005:src0_endofpacket -> ddr2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_005_src0_valid;                                                                      // cmd_xbar_demux_005:src0_valid -> ddr2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_005_src0_startofpacket;                                                              // cmd_xbar_demux_005:src0_startofpacket -> ddr2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [94:0] cmd_xbar_demux_005_src0_data;                                                                       // cmd_xbar_demux_005:src0_data -> ddr2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [0:0] cmd_xbar_demux_005_src0_channel;                                                                    // cmd_xbar_demux_005:src0_channel -> ddr2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_030_src0_endofpacket;                                                                // rsp_xbar_demux_030:src0_endofpacket -> cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_030_src0_valid;                                                                      // rsp_xbar_demux_030:src0_valid -> cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_030_src0_startofpacket;                                                              // rsp_xbar_demux_030:src0_startofpacket -> cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [94:0] rsp_xbar_demux_030_src0_data;                                                                       // rsp_xbar_demux_030:src0_data -> cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [0:0] rsp_xbar_demux_030_src0_channel;                                                                    // rsp_xbar_demux_030:src0_channel -> cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          addr_router_005_src_endofpacket;                                                                    // addr_router_005:src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire          addr_router_005_src_valid;                                                                          // addr_router_005:src_valid -> cmd_xbar_demux_005:sink_valid
	wire          addr_router_005_src_startofpacket;                                                                  // addr_router_005:src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire   [94:0] addr_router_005_src_data;                                                                           // addr_router_005:src_data -> cmd_xbar_demux_005:sink_data
	wire    [0:0] addr_router_005_src_channel;                                                                        // addr_router_005:src_channel -> cmd_xbar_demux_005:sink_channel
	wire          addr_router_005_src_ready;                                                                          // cmd_xbar_demux_005:sink_ready -> addr_router_005:src_ready
	wire          rsp_xbar_demux_030_src0_ready;                                                                      // cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_030:src0_ready
	wire          cmd_xbar_demux_005_src0_ready;                                                                      // ddr2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_005:src0_ready
	wire          id_router_030_src_endofpacket;                                                                      // id_router_030:src_endofpacket -> rsp_xbar_demux_030:sink_endofpacket
	wire          id_router_030_src_valid;                                                                            // id_router_030:src_valid -> rsp_xbar_demux_030:sink_valid
	wire          id_router_030_src_startofpacket;                                                                    // id_router_030:src_startofpacket -> rsp_xbar_demux_030:sink_startofpacket
	wire   [94:0] id_router_030_src_data;                                                                             // id_router_030:src_data -> rsp_xbar_demux_030:sink_data
	wire    [0:0] id_router_030_src_channel;                                                                          // id_router_030:src_channel -> rsp_xbar_demux_030:sink_channel
	wire          id_router_030_src_ready;                                                                            // rsp_xbar_demux_030:sink_ready -> id_router_030:src_ready
	wire          crosser_out_endofpacket;                                                                            // crosser:out_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_out_valid;                                                                                  // crosser:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_out_startofpacket;                                                                          // crosser:out_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] crosser_out_data;                                                                                   // crosser:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [23:0] crosser_out_channel;                                                                                // crosser:out_channel -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                // cmd_xbar_demux_003:src0_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                      // cmd_xbar_demux_003:src0_valid -> crosser:in_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                              // cmd_xbar_demux_003:src0_startofpacket -> crosser:in_startofpacket
	wire   [84:0] cmd_xbar_demux_003_src0_data;                                                                       // cmd_xbar_demux_003:src0_data -> crosser:in_data
	wire   [23:0] cmd_xbar_demux_003_src0_channel;                                                                    // cmd_xbar_demux_003:src0_channel -> crosser:in_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                      // crosser:in_ready -> cmd_xbar_demux_003:src0_ready
	wire          crosser_001_out_endofpacket;                                                                        // crosser_001:out_endofpacket -> cmd_xbar_mux_021:sink1_endofpacket
	wire          crosser_001_out_valid;                                                                              // crosser_001:out_valid -> cmd_xbar_mux_021:sink1_valid
	wire          crosser_001_out_startofpacket;                                                                      // crosser_001:out_startofpacket -> cmd_xbar_mux_021:sink1_startofpacket
	wire   [84:0] crosser_001_out_data;                                                                               // crosser_001:out_data -> cmd_xbar_mux_021:sink1_data
	wire   [23:0] crosser_001_out_channel;                                                                            // crosser_001:out_channel -> cmd_xbar_mux_021:sink1_channel
	wire          crosser_001_out_ready;                                                                              // cmd_xbar_mux_021:sink1_ready -> crosser_001:out_ready
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                                // cmd_xbar_demux_004:src0_endofpacket -> crosser_001:in_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                      // cmd_xbar_demux_004:src0_valid -> crosser_001:in_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                              // cmd_xbar_demux_004:src0_startofpacket -> crosser_001:in_startofpacket
	wire   [84:0] cmd_xbar_demux_004_src0_data;                                                                       // cmd_xbar_demux_004:src0_data -> crosser_001:in_data
	wire   [23:0] cmd_xbar_demux_004_src0_channel;                                                                    // cmd_xbar_demux_004:src0_channel -> crosser_001:in_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                      // crosser_001:in_ready -> cmd_xbar_demux_004:src0_ready
	wire          crosser_002_out_endofpacket;                                                                        // crosser_002:out_endofpacket -> cmd_xbar_mux_022:sink1_endofpacket
	wire          crosser_002_out_valid;                                                                              // crosser_002:out_valid -> cmd_xbar_mux_022:sink1_valid
	wire          crosser_002_out_startofpacket;                                                                      // crosser_002:out_startofpacket -> cmd_xbar_mux_022:sink1_startofpacket
	wire   [84:0] crosser_002_out_data;                                                                               // crosser_002:out_data -> cmd_xbar_mux_022:sink1_data
	wire   [23:0] crosser_002_out_channel;                                                                            // crosser_002:out_channel -> cmd_xbar_mux_022:sink1_channel
	wire          crosser_002_out_ready;                                                                              // cmd_xbar_mux_022:sink1_ready -> crosser_002:out_ready
	wire          cmd_xbar_demux_004_src1_endofpacket;                                                                // cmd_xbar_demux_004:src1_endofpacket -> crosser_002:in_endofpacket
	wire          cmd_xbar_demux_004_src1_valid;                                                                      // cmd_xbar_demux_004:src1_valid -> crosser_002:in_valid
	wire          cmd_xbar_demux_004_src1_startofpacket;                                                              // cmd_xbar_demux_004:src1_startofpacket -> crosser_002:in_startofpacket
	wire   [84:0] cmd_xbar_demux_004_src1_data;                                                                       // cmd_xbar_demux_004:src1_data -> crosser_002:in_data
	wire   [23:0] cmd_xbar_demux_004_src1_channel;                                                                    // cmd_xbar_demux_004:src1_channel -> crosser_002:in_channel
	wire          cmd_xbar_demux_004_src1_ready;                                                                      // crosser_002:in_ready -> cmd_xbar_demux_004:src1_ready
	wire          crosser_003_out_endofpacket;                                                                        // crosser_003:out_endofpacket -> rsp_xbar_mux_003:sink0_endofpacket
	wire          crosser_003_out_valid;                                                                              // crosser_003:out_valid -> rsp_xbar_mux_003:sink0_valid
	wire          crosser_003_out_startofpacket;                                                                      // crosser_003:out_startofpacket -> rsp_xbar_mux_003:sink0_startofpacket
	wire   [84:0] crosser_003_out_data;                                                                               // crosser_003:out_data -> rsp_xbar_mux_003:sink0_data
	wire   [23:0] crosser_003_out_channel;                                                                            // crosser_003:out_channel -> rsp_xbar_mux_003:sink0_channel
	wire          crosser_003_out_ready;                                                                              // rsp_xbar_mux_003:sink0_ready -> crosser_003:out_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                // rsp_xbar_demux_006:src0_endofpacket -> crosser_003:in_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                      // rsp_xbar_demux_006:src0_valid -> crosser_003:in_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                              // rsp_xbar_demux_006:src0_startofpacket -> crosser_003:in_startofpacket
	wire   [84:0] rsp_xbar_demux_006_src0_data;                                                                       // rsp_xbar_demux_006:src0_data -> crosser_003:in_data
	wire   [23:0] rsp_xbar_demux_006_src0_channel;                                                                    // rsp_xbar_demux_006:src0_channel -> crosser_003:in_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                      // crosser_003:in_ready -> rsp_xbar_demux_006:src0_ready
	wire          crosser_004_out_endofpacket;                                                                        // crosser_004:out_endofpacket -> rsp_xbar_mux_004:sink0_endofpacket
	wire          crosser_004_out_valid;                                                                              // crosser_004:out_valid -> rsp_xbar_mux_004:sink0_valid
	wire          crosser_004_out_startofpacket;                                                                      // crosser_004:out_startofpacket -> rsp_xbar_mux_004:sink0_startofpacket
	wire   [84:0] crosser_004_out_data;                                                                               // crosser_004:out_data -> rsp_xbar_mux_004:sink0_data
	wire   [23:0] crosser_004_out_channel;                                                                            // crosser_004:out_channel -> rsp_xbar_mux_004:sink0_channel
	wire          crosser_004_out_ready;                                                                              // rsp_xbar_mux_004:sink0_ready -> crosser_004:out_ready
	wire          rsp_xbar_demux_021_src1_endofpacket;                                                                // rsp_xbar_demux_021:src1_endofpacket -> crosser_004:in_endofpacket
	wire          rsp_xbar_demux_021_src1_valid;                                                                      // rsp_xbar_demux_021:src1_valid -> crosser_004:in_valid
	wire          rsp_xbar_demux_021_src1_startofpacket;                                                              // rsp_xbar_demux_021:src1_startofpacket -> crosser_004:in_startofpacket
	wire   [84:0] rsp_xbar_demux_021_src1_data;                                                                       // rsp_xbar_demux_021:src1_data -> crosser_004:in_data
	wire   [23:0] rsp_xbar_demux_021_src1_channel;                                                                    // rsp_xbar_demux_021:src1_channel -> crosser_004:in_channel
	wire          rsp_xbar_demux_021_src1_ready;                                                                      // crosser_004:in_ready -> rsp_xbar_demux_021:src1_ready
	wire          crosser_005_out_endofpacket;                                                                        // crosser_005:out_endofpacket -> rsp_xbar_mux_004:sink1_endofpacket
	wire          crosser_005_out_valid;                                                                              // crosser_005:out_valid -> rsp_xbar_mux_004:sink1_valid
	wire          crosser_005_out_startofpacket;                                                                      // crosser_005:out_startofpacket -> rsp_xbar_mux_004:sink1_startofpacket
	wire   [84:0] crosser_005_out_data;                                                                               // crosser_005:out_data -> rsp_xbar_mux_004:sink1_data
	wire   [23:0] crosser_005_out_channel;                                                                            // crosser_005:out_channel -> rsp_xbar_mux_004:sink1_channel
	wire          crosser_005_out_ready;                                                                              // rsp_xbar_mux_004:sink1_ready -> crosser_005:out_ready
	wire          rsp_xbar_demux_022_src1_endofpacket;                                                                // rsp_xbar_demux_022:src1_endofpacket -> crosser_005:in_endofpacket
	wire          rsp_xbar_demux_022_src1_valid;                                                                      // rsp_xbar_demux_022:src1_valid -> crosser_005:in_valid
	wire          rsp_xbar_demux_022_src1_startofpacket;                                                              // rsp_xbar_demux_022:src1_startofpacket -> crosser_005:in_startofpacket
	wire   [84:0] rsp_xbar_demux_022_src1_data;                                                                       // rsp_xbar_demux_022:src1_data -> crosser_005:in_data
	wire   [23:0] rsp_xbar_demux_022_src1_channel;                                                                    // rsp_xbar_demux_022:src1_channel -> crosser_005:in_channel
	wire          rsp_xbar_demux_022_src1_ready;                                                                      // crosser_005:in_ready -> rsp_xbar_demux_022:src1_ready
	wire    [5:0] limiter_cmd_valid_data;                                                                             // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [23:0] limiter_001_cmd_valid_data;                                                                         // limiter_001:cmd_src_valid -> cmd_xbar_demux_003:sink_valid
	wire          irq_mapper_receiver5_irq;                                                                           // epcs_flash:irq -> irq_mapper:receiver5_irq
	wire          irq_mapper_receiver6_irq;                                                                           // dma_0:dma_ctl_irq -> irq_mapper:receiver6_irq
	wire   [31:0] nios2_d_irq_irq;                                                                                    // irq_mapper:sender_irq -> nios2:d_irq
	wire          irq_mapper_receiver0_irq;                                                                           // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                                                      // jtag_uart_0:av_irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver1_irq;                                                                           // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                                                                  // systimer:irq -> irq_synchronizer_001:receiver_irq
	wire          irq_mapper_receiver2_irq;                                                                           // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire    [0:0] irq_synchronizer_002_receiver_irq;                                                                  // pio_key:irq -> irq_synchronizer_002:receiver_irq
	wire          irq_mapper_receiver3_irq;                                                                           // irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	wire    [0:0] irq_synchronizer_003_receiver_irq;                                                                  // uart_0:irq -> irq_synchronizer_003:receiver_irq
	wire          irq_mapper_receiver4_irq;                                                                           // irq_synchronizer_004:sender_irq -> irq_mapper:receiver4_irq
	wire    [0:0] irq_synchronizer_004_receiver_irq;                                                                  // spi_0:irq -> irq_synchronizer_004:receiver_irq
	wire          irq_mapper_receiver7_irq;                                                                           // irq_synchronizer_005:sender_irq -> irq_mapper:receiver7_irq
	wire    [0:0] irq_synchronizer_005_receiver_irq;                                                                  // timestamp:irq -> irq_synchronizer_005:receiver_irq
	wire          irq_mapper_receiver8_irq;                                                                           // irq_synchronizer_006:sender_irq -> irq_mapper:receiver8_irq
	wire    [0:0] irq_synchronizer_006_receiver_irq;                                                                  // spi_ad5781:irq -> irq_synchronizer_006:receiver_irq
	wire          irq_mapper_receiver9_irq;                                                                           // irq_synchronizer_007:sender_irq -> irq_mapper:receiver9_irq
	wire    [0:0] irq_synchronizer_007_receiver_irq;                                                                  // oc_i2c_master_0:wb_inta_o -> irq_synchronizer_007:receiver_irq
	wire          irq_mapper_receiver10_irq;                                                                          // irq_synchronizer_008:sender_irq -> irq_mapper:receiver10_irq
	wire    [0:0] irq_synchronizer_008_receiver_irq;                                                                  // spi_master_0:interrupt -> irq_synchronizer_008:receiver_irq
	wire          irq_mapper_receiver11_irq;                                                                          // irq_synchronizer_009:sender_irq -> irq_mapper:receiver11_irq
	wire    [0:0] irq_synchronizer_009_receiver_irq;                                                                  // ad9266:irq -> irq_synchronizer_009:receiver_irq

	nios2_nios2 nios2 (
		.clk                                   (nios_clk_clk),                                                       //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                    //                   reset_n.reset_n
		.d_address                             (nios2_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2_data_master_read),                                             //                          .read
		.d_readdata                            (nios2_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2_data_master_write),                                            //                          .write
		.d_writedata                           (nios2_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2_instruction_master_waitrequest),                               //                          .waitrequest
		.i_readdatavalid                       (nios2_instruction_master_readdatavalid),                             //                          .readdatavalid
		.d_irq                                 (nios2_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	nios2_onchip_ram onchip_ram (
		.clk        (nios_clk_clk),                                            //   clk1.clk
		.address    (onchip_ram_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_ram_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_ram_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_ram_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_ram_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_ram_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_ram_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                           // reset1.reset
	);

	nios2_sysid sysid (
		.clock    (altpll_0_c0_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                         //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	nios2_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c0_clk),                                                          //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_receiver_irq)                                             //               irq.irq
	);

	nios2_ddr2 ddr2 (
		.local_address        (ddr2_s1_translator_avalon_anti_slave_0_address),            //                  s1.address
		.local_write_req      (ddr2_s1_translator_avalon_anti_slave_0_write),              //                    .write
		.local_read_req       (ddr2_s1_translator_avalon_anti_slave_0_read),               //                    .read
		.local_burstbegin     (ddr2_s1_translator_avalon_anti_slave_0_beginbursttransfer), //                    .beginbursttransfer
		.local_ready          (ddr2_s1_translator_avalon_anti_slave_0_waitrequest),        //                    .waitrequest_n
		.local_rdata          (ddr2_s1_translator_avalon_anti_slave_0_readdata),           //                    .readdata
		.local_rdata_valid    (ddr2_s1_translator_avalon_anti_slave_0_readdatavalid),      //                    .readdatavalid
		.local_wdata          (ddr2_s1_translator_avalon_anti_slave_0_writedata),          //                    .writedata
		.local_be             (ddr2_s1_translator_avalon_anti_slave_0_byteenable),         //                    .byteenable
		.local_size           (ddr2_s1_translator_avalon_anti_slave_0_burstcount),         //                    .burstcount
		.local_refresh_ack    (),                                                          // external_connection.export
		.local_init_done      (),                                                          //                    .export
		.reset_phy_clk_n      (),                                                          //                    .export
		.local_self_rfsh_req  (),                                                          //                    .export
		.local_self_rfsh_chip (),                                                          //                    .export
		.local_self_rfsh_ack  (),                                                          //                    .export
		.mem_odt              (ddr2_mem_odt),                                              //              memory.mem_odt
		.mem_clk              (ddr2_mem_clk),                                              //                    .mem_clk
		.mem_clk_n            (ddr2_mem_clk_n),                                            //                    .mem_clk_n
		.mem_cs_n             (ddr2_mem_cs_n),                                             //                    .mem_cs_n
		.mem_cke              (ddr2_mem_cke),                                              //                    .mem_cke
		.mem_addr             (ddr2_mem_addr),                                             //                    .mem_addr
		.mem_ba               (ddr2_mem_ba),                                               //                    .mem_ba
		.mem_ras_n            (ddr2_mem_ras_n),                                            //                    .mem_ras_n
		.mem_cas_n            (ddr2_mem_cas_n),                                            //                    .mem_cas_n
		.mem_we_n             (ddr2_mem_we_n),                                             //                    .mem_we_n
		.mem_dq               (ddr2_mem_dq),                                               //                    .mem_dq
		.mem_dqs              (ddr2_mem_dqs),                                              //                    .mem_dqs
		.mem_dm               (ddr2_mem_dm),                                               //                    .mem_dm
		.pll_ref_clk          (altpll_0_c1_clk),                                           //              refclk.clk
		.soft_reset_n         (~rst_controller_002_reset_out_reset),                       //        soft_reset_n.reset_n
		.global_reset_n       (~rst_controller_003_reset_out_reset),                       //      global_reset_n.reset_n
		.reset_request_n      (ddr2_reset_request_n_reset),                                //     reset_request_n.reset_n
		.phy_clk              (ddr2_sysclk_clk),                                           //              sysclk.clk
		.aux_full_rate_clk    (),                                                          //             auxfull.clk
		.aux_half_rate_clk    ()                                                           //             auxhalf.clk
	);

	nios2_systimer systimer (
		.clk        (altpll_0_c0_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                   // reset.reset_n
		.address    (systimer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (systimer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (systimer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (systimer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~systimer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)                      //   irq.irq
	);

	nios2_pio_led pio_led (
		.clk        (altpll_0_c0_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address    (pio_led_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_led_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_led_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_led_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_led_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_export)                                            // external_connection.export
	);

	nios2_pio_key pio_key (
		.clk        (altpll_0_c0_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address    (pio_key_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_key_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_key_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_key_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_key_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (key_export),                                           // external_connection.export
		.irq        (irq_synchronizer_002_receiver_irq)                     //                 irq.irq
	);

	nios2_uart_0 uart_0 (
		.clk           (altpll_0_c0_clk),                                        //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address       (uart_0_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (uart_0_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (uart_0_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~uart_0_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~uart_0_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (uart_0_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (uart_0_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                       //                    .dataavailable
		.readyfordata  (),                                                       //                    .readyfordata
		.rxd           (uart_rxd),                                               // external_connection.export
		.txd           (uart_txd),                                               //                    .export
		.irq           (irq_synchronizer_003_receiver_irq)                       //                 irq.irq
	);

	nios2_spi_0 spi_0 (
		.clk           (altpll_0_c0_clk),                                                  //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                              //            reset.reset_n
		.data_from_cpu (spi_0_spi_control_port_translator_avalon_anti_slave_0_writedata),  // spi_control_port.writedata
		.data_to_cpu   (spi_0_spi_control_port_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.mem_addr      (spi_0_spi_control_port_translator_avalon_anti_slave_0_address),    //                 .address
		.read_n        (~spi_0_spi_control_port_translator_avalon_anti_slave_0_read),      //                 .read_n
		.spi_select    (spi_0_spi_control_port_translator_avalon_anti_slave_0_chipselect), //                 .chipselect
		.write_n       (~spi_0_spi_control_port_translator_avalon_anti_slave_0_write),     //                 .write_n
		.irq           (irq_synchronizer_004_receiver_irq),                                //              irq.irq
		.MISO          (spi_dp_MISO),                                                      //         external.export
		.MOSI          (spi_dp_MOSI),                                                      //                 .export
		.SCLK          (spi_dp_SCLK),                                                      //                 .export
		.SS_n          (spi_dp_SS_n)                                                       //                 .export
	);

	nios2_epcs_flash epcs_flash (
		.clk           (nios_clk_clk),                                                           //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.address       (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_address),    // epcs_control_port.address
		.chipselect    (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_chipselect), //                  .chipselect
		.dataavailable (),                                                                       //                  .dataavailable
		.endofpacket   (),                                                                       //                  .endofpacket
		.read_n        (~epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_read),      //                  .read_n
		.readdata      (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_readdata),   //                  .readdata
		.readyfordata  (),                                                                       //                  .readyfordata
		.write_n       (~epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_write),     //                  .write_n
		.writedata     (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver5_irq),                                               //               irq.irq
		.dclk          (epcs_flash_dclk),                                                        //          external.export
		.sce           (epcs_flash_sce),                                                         //                  .export
		.sdo           (epcs_flash_sdo),                                                         //                  .export
		.data0         (epcs_flash_data0)                                                        //                  .export
	);

	nios2_altpll_0 altpll_0 (
		.clk       (clk_clk),                                                     //       inclk_interface.clk
		.reset     (rst_controller_004_reset_out_reset),                          // inclk_interface_reset.reset
		.read      (altpll_0_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (altpll_0_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (altpll_0_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (altpll_0_c0_clk),                                             //                    c0.clk
		.c1        (altpll_0_c1_clk),                                             //                    c1.clk
		.c2        (nios_clk_clk),                                                //                    c2.clk
		.c3        (),                                                            //            c3_conduit.export
		.areset    (),                                                            //        areset_conduit.export
		.locked    (),                                                            //        locked_conduit.export
		.phasedone ()                                                             //     phasedone_conduit.export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (16),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) slow_peripheral_bridge (
		.m0_clk           (altpll_0_c0_clk),                                                        //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                                     // m0_reset.reset
		.s0_clk           (nios_clk_clk),                                                           //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                                         // s0_reset.reset
		.s0_waitrequest   (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (slow_peripheral_bridge_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (slow_peripheral_bridge_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (slow_peripheral_bridge_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (slow_peripheral_bridge_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (slow_peripheral_bridge_m0_writedata),                                    //         .writedata
		.m0_address       (slow_peripheral_bridge_m0_address),                                      //         .address
		.m0_write         (slow_peripheral_bridge_m0_write),                                        //         .write
		.m0_read          (slow_peripheral_bridge_m0_read),                                         //         .read
		.m0_byteenable    (slow_peripheral_bridge_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (slow_peripheral_bridge_m0_debugaccess)                                   //         .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (26),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) cpu_ddr2_clock_bridge (
		.m0_clk           (ddr2_sysclk_clk),                                                       //   m0_clk.clk
		.m0_reset         (rst_controller_005_reset_out_reset),                                    // m0_reset.reset
		.s0_clk           (nios_clk_clk),                                                          //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                                        // s0_reset.reset
		.s0_waitrequest   (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (cpu_ddr2_clock_bridge_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (cpu_ddr2_clock_bridge_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (cpu_ddr2_clock_bridge_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (cpu_ddr2_clock_bridge_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (cpu_ddr2_clock_bridge_m0_writedata),                                    //         .writedata
		.m0_address       (cpu_ddr2_clock_bridge_m0_address),                                      //         .address
		.m0_write         (cpu_ddr2_clock_bridge_m0_write),                                        //         .write
		.m0_read          (cpu_ddr2_clock_bridge_m0_read),                                         //         .read
		.m0_byteenable    (cpu_ddr2_clock_bridge_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (cpu_ddr2_clock_bridge_m0_debugaccess)                                   //         .debugaccess
	);

	nios2_dma_0 dma_0 (
		.clk                (nios_clk_clk),                                                       //                clk.clk
		.system_reset_n     (~rst_controller_reset_out_reset),                                    //              reset.reset_n
		.dma_ctl_address    (dma_0_control_port_slave_translator_avalon_anti_slave_0_address),    // control_port_slave.address
		.dma_ctl_chipselect (dma_0_control_port_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.dma_ctl_readdata   (dma_0_control_port_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.dma_ctl_write_n    (~dma_0_control_port_slave_translator_avalon_anti_slave_0_write),     //                   .write_n
		.dma_ctl_writedata  (dma_0_control_port_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_receiver6_irq),                                           //                irq.irq
		.read_address       (dma_0_read_master_address),                                          //        read_master.address
		.read_chipselect    (dma_0_read_master_chipselect),                                       //                   .chipselect
		.read_read_n        (dma_0_read_master_read),                                             //                   .read_n
		.read_readdata      (dma_0_read_master_readdata),                                         //                   .readdata
		.read_readdatavalid (dma_0_read_master_readdatavalid),                                    //                   .readdatavalid
		.read_waitrequest   (dma_0_read_master_waitrequest),                                      //                   .waitrequest
		.write_address      (dma_0_write_master_address),                                         //       write_master.address
		.write_chipselect   (dma_0_write_master_chipselect),                                      //                   .chipselect
		.write_waitrequest  (dma_0_write_master_waitrequest),                                     //                   .waitrequest
		.write_write_n      (dma_0_write_master_write),                                           //                   .write_n
		.write_writedata    (dma_0_write_master_writedata),                                       //                   .writedata
		.write_byteenable   (dma_0_write_master_byteenable)                                       //                   .byteenable
	);

	nios2_timestamp timestamp (
		.clk        (altpll_0_c0_clk),                                        //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    // reset.reset_n
		.address    (timestamp_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timestamp_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timestamp_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timestamp_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timestamp_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_005_receiver_irq)                       //   irq.irq
	);

	nios2_spi_ad5781 spi_ad5781 (
		.clk           (altpll_0_c0_clk),                                                       //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                                   //            reset.reset_n
		.data_from_cpu (spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_writedata),  // spi_control_port.writedata
		.data_to_cpu   (spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.mem_addr      (spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_address),    //                 .address
		.read_n        (~spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_read),      //                 .read_n
		.spi_select    (spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_chipselect), //                 .chipselect
		.write_n       (~spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_write),     //                 .write_n
		.irq           (irq_synchronizer_006_receiver_irq),                                     //              irq.irq
		.MISO          (spi_ad5781_MISO),                                                       //         external.export
		.MOSI          (spi_ad5781_MOSI),                                                       //                 .export
		.SCLK          (spi_ad5781_SCLK),                                                       //                 .export
		.SS_n          (spi_ad5781_SS_n)                                                        //                 .export
	);

	ad9245 ad9245_2 (
		.clk        (altpll_0_c0_clk),                                       //     clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                   //   reset.reset_n
		.chipselect (ad9245_2_s1_translator_avalon_anti_slave_0_chipselect), //      s1.chipselect
		.read       (ad9245_2_s1_translator_avalon_anti_slave_0_read),       //        .read
		.readdata   (ad9245_2_s1_translator_avalon_anti_slave_0_readdata),   //        .readdata
		.ad_data    (ad9245_2_ad_data_export)                                // ad_data.export
	);

	ad9245 ad9245_1 (
		.clk        (altpll_0_c0_clk),                                       //     clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                   //   reset.reset_n
		.chipselect (ad9245_1_s1_translator_avalon_anti_slave_0_chipselect), //      s1.chipselect
		.read       (ad9245_1_s1_translator_avalon_anti_slave_0_read),       //        .read
		.readdata   (ad9245_1_s1_translator_avalon_anti_slave_0_readdata),   //        .readdata
		.ad_data    (ad9245_1_ad_data_export)                                // ad_data.export
	);

	clk_gen #(
		.clk_num (8)
	) clk_gen (
		.reset_n    (~rst_controller_001_reset_out_reset),                  //      reset.reset_n
		.chipselect (clk_gen_s1_translator_avalon_anti_slave_0_chipselect), //         s1.chipselect
		.address    (clk_gen_s1_translator_avalon_anti_slave_0_address),    //           .address
		.read       (clk_gen_s1_translator_avalon_anti_slave_0_read),       //           .read
		.write      (clk_gen_s1_translator_avalon_anti_slave_0_write),      //           .write
		.readdata   (clk_gen_s1_translator_avalon_anti_slave_0_readdata),   //           .readdata
		.writedata  (clk_gen_s1_translator_avalon_anti_slave_0_writedata),  //           .writedata
		.clk        (altpll_0_c0_clk),                                      //        clk.clk
		.clk_source (nios_clk_clk),                                         // clk_source.clk
		.clk_out    (clk_gen_clk_out_export)                                //    clk_out.export
	);

	oc_i2c_master oc_i2c_master_0 (
		.wb_clk_i   (altpll_0_c0_clk),                                                 //       s1_clk.clk
		.wb_rst_i   (rst_controller_001_reset_out_reset),                              // s1_clk_reset.reset
		.wb_ack_o   (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_waitrequest),   //           s1.waitrequest_n
		.wb_adr_i   (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_address),       //             .address
		.wb_dat_i   (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_writedata),     //             .writedata
		.wb_dat_o   (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_readdata),      //             .readdata
		.wb_stb_i   (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_begintransfer), //             .begintransfer
		.wb_we_i    (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_write),         //             .write
		.wb_cyc_i   (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_chipselect),    //             .chipselect
		.scl_pad_io (oc_i2c_master_scl_pad_io),                                        //       global.export
		.sda_pad_io (oc_i2c_master_sda_pad_io),                                        //             .export
		.wb_inta_o  (irq_synchronizer_007_receiver_irq)                                //       s1_irq.irq
	);

	spi_master #(
		.numberOfSlaves (1),
		.clk_pol        (1),
		.clk_pha        (0)
	) spi_master_0 (
		.clk        (altpll_0_c0_clk),                                           //       clock.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                       //       reset.reset_n
		.miso       (spi_master_miso),                                           // conduit_end.export
		.mosi       (spi_master_mosi),                                           //            .export
		.sclk       (spi_master_sclk),                                           //            .export
		.ss         (spi_master_ss),                                             //            .export
		.chipselect (spi_master_0_s1_translator_avalon_anti_slave_0_chipselect), //          s1.chipselect
		.address    (spi_master_0_s1_translator_avalon_anti_slave_0_address),    //            .address
		.read       (spi_master_0_s1_translator_avalon_anti_slave_0_read),       //            .read
		.write      (spi_master_0_s1_translator_avalon_anti_slave_0_write),      //            .write
		.readdata   (spi_master_0_s1_translator_avalon_anti_slave_0_readdata),   //            .readdata
		.writedata  (spi_master_0_s1_translator_avalon_anti_slave_0_writedata),  //            .writedata
		.interrupt  (irq_synchronizer_008_receiver_irq)                          //   interrupt.irq
	);

	nios2_ad9266 ad9266 (
		.clk           (altpll_0_c0_clk),                                                   //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                               //            reset.reset_n
		.data_from_cpu (ad9266_spi_control_port_translator_avalon_anti_slave_0_writedata),  // spi_control_port.writedata
		.data_to_cpu   (ad9266_spi_control_port_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.mem_addr      (ad9266_spi_control_port_translator_avalon_anti_slave_0_address),    //                 .address
		.read_n        (~ad9266_spi_control_port_translator_avalon_anti_slave_0_read),      //                 .read_n
		.spi_select    (ad9266_spi_control_port_translator_avalon_anti_slave_0_chipselect), //                 .chipselect
		.write_n       (~ad9266_spi_control_port_translator_avalon_anti_slave_0_write),     //                 .write_n
		.irq           (irq_synchronizer_009_receiver_irq),                                 //              irq.irq
		.MISO          (ad9266_MISO),                                                       //         external.export
		.MOSI          (ad9266_MOSI),                                                       //                 .export
		.SCLK          (ad9266_SCLK),                                                       //                 .export
		.SS_n          (ad9266_SS_n)                                                        //                 .export
	);

	dac2904 dac2904_1 (
		.reset_n            (~rst_controller_001_reset_out_reset),                     //      reset.reset_n
		.clk                (altpll_0_c0_clk),                                         //        clk.clk
		.dac_data           (dac2904_1_dac_data_export),                               //   dac_data.export
		.avs_s0_chipselect  (dac2904_1_s0_translator_avalon_anti_slave_0_chipselect),  //         s0.chipselect
		.avs_s0_write       (dac2904_1_s0_translator_avalon_anti_slave_0_write),       //           .write
		.avs_s0_writedata   (dac2904_1_s0_translator_avalon_anti_slave_0_writedata),   //           .writedata
		.avs_s0_waitrequest (dac2904_1_s0_translator_avalon_anti_slave_0_waitrequest), //           .waitrequest
		.sample_clock       (dac2904_1_sample_clk_clk)                                 // sample_clk.clk
	);

	dac2904 dac2904_2 (
		.reset_n            (~rst_controller_001_reset_out_reset),                     //      reset.reset_n
		.clk                (altpll_0_c0_clk),                                         //        clk.clk
		.dac_data           (dac2904_2_dac_data_export),                               //   dac_data.export
		.avs_s0_chipselect  (dac2904_2_s0_translator_avalon_anti_slave_0_chipselect),  //         s0.chipselect
		.avs_s0_write       (dac2904_2_s0_translator_avalon_anti_slave_0_write),       //           .write
		.avs_s0_writedata   (dac2904_2_s0_translator_avalon_anti_slave_0_writedata),   //           .writedata
		.avs_s0_waitrequest (dac2904_2_s0_translator_avalon_anti_slave_0_waitrequest), //           .waitrequest
		.sample_clock       (dac2904_2_sample_clk_clk)                                 // sample_clk.clk
	);

	dac2904 dac2904_3 (
		.reset_n            (~rst_controller_001_reset_out_reset),                     //      reset.reset_n
		.clk                (altpll_0_c0_clk),                                         //        clk.clk
		.dac_data           (dac2904_3_dac_data_export),                               //   dac_data.export
		.avs_s0_chipselect  (dac2904_3_s0_translator_avalon_anti_slave_0_chipselect),  //         s0.chipselect
		.avs_s0_write       (dac2904_3_s0_translator_avalon_anti_slave_0_write),       //           .write
		.avs_s0_writedata   (dac2904_3_s0_translator_avalon_anti_slave_0_writedata),   //           .writedata
		.avs_s0_waitrequest (dac2904_3_s0_translator_avalon_anti_slave_0_waitrequest), //           .waitrequest
		.sample_clock       (dac2904_3_sample_clk_clk)                                 // sample_clk.clk
	);

	dac2904 dac2904_4 (
		.reset_n            (~rst_controller_001_reset_out_reset),                     //      reset.reset_n
		.clk                (altpll_0_c0_clk),                                         //        clk.clk
		.dac_data           (dac2904_4_dac_data_export),                               //   dac_data.export
		.avs_s0_chipselect  (dac2904_4_s0_translator_avalon_anti_slave_0_chipselect),  //         s0.chipselect
		.avs_s0_write       (dac2904_4_s0_translator_avalon_anti_slave_0_write),       //           .write
		.avs_s0_writedata   (dac2904_4_s0_translator_avalon_anti_slave_0_writedata),   //           .writedata
		.avs_s0_waitrequest (dac2904_4_s0_translator_avalon_anti_slave_0_waitrequest), //           .waitrequest
		.sample_clock       (dac2904_4_sample_clk_clk)                                 // sample_clk.clk
	);

	wave_gen #(
		.AmpMax       (14'b11111111111111),
		.AmpMin       (14'b00000000000000),
		.FreqDiv      (34'b0000000000000000000000000000010100),
		.SamplePonint (13'b0000100000000)
	) wave_gen_0 (
		.clk               (altpll_0_c0_clk),                                         //      clock.clk
		.reset_n           (~rst_controller_001_reset_out_reset),                     //      reset.reset_n
		.avs_s0_chipselect (wave_gen_0_s0_translator_avalon_anti_slave_0_chipselect), //         s0.chipselect
		.avs_s0_write      (wave_gen_0_s0_translator_avalon_anti_slave_0_write),      //           .write
		.avs_s0_read       (wave_gen_0_s0_translator_avalon_anti_slave_0_read),       //           .read
		.avs_s0_writedata  (wave_gen_0_s0_translator_avalon_anti_slave_0_writedata),  //           .writedata
		.avs_s0_readdata   (wave_gen_0_s0_translator_avalon_anti_slave_0_readdata),   //           .readdata
		.avs_s0_address    (wave_gen_0_s0_translator_avalon_anti_slave_0_address),    //           .address
		.clk_source        (nios_clk_clk),                                            // clk_source.clk
		.dac               (wave_gen_0_dac_export)                                    //        dac.export
	);

	demodulation #(
		.Sample1Start (18'b000000000000100000),
		.Sample2Start (18'b000000000010000000),
		.Sample1Num   (18'b000000000000100000),
		.Sample2Num   (18'b000000000000100000),
		.FreqDiv      (34'b0000000000000000000000000000000001)
	) demodulation_0 (
		.clk               (altpll_0_c0_clk),                                             //      clock.clk
		.reset_n           (~rst_controller_001_reset_out_reset),                         //      reset.reset_n
		.avs_s0_chipselect (demodulation_0_s0_translator_avalon_anti_slave_0_chipselect), //         s0.chipselect
		.avs_s0_write      (demodulation_0_s0_translator_avalon_anti_slave_0_write),      //           .write
		.avs_s0_read       (demodulation_0_s0_translator_avalon_anti_slave_0_read),       //           .read
		.avs_s0_writedata  (demodulation_0_s0_translator_avalon_anti_slave_0_writedata),  //           .writedata
		.avs_s0_readdata   (demodulation_0_s0_translator_avalon_anti_slave_0_readdata),   //           .readdata
		.avs_s0_address    (demodulation_0_s0_translator_avalon_anti_slave_0_address),    //           .address
		.clk_source        (nios_clk_clk),                                                // clk_source.clk
		.dac               (demodulation_0_ad_da_dac),                                    //      ad_da.export
		.ad                (demodulation_0_ad_da_ad),                                     //           .export
		.modulation_wave   (demodulation_0_ad_da_modulation_wave)                         //           .export
	);

	wave_gen #(
		.AmpMax       (14'b11111111111111),
		.AmpMin       (14'b00000000000000),
		.FreqDiv      (34'b0000000000000000000000000000010100),
		.SamplePonint (13'b0000100000000)
	) wave_gen_1 (
		.clk               (altpll_0_c0_clk),                                         //      clock.clk
		.reset_n           (~rst_controller_001_reset_out_reset),                     //      reset.reset_n
		.avs_s0_chipselect (wave_gen_1_s0_translator_avalon_anti_slave_0_chipselect), //         s0.chipselect
		.avs_s0_write      (wave_gen_1_s0_translator_avalon_anti_slave_0_write),      //           .write
		.avs_s0_read       (wave_gen_1_s0_translator_avalon_anti_slave_0_read),       //           .read
		.avs_s0_writedata  (wave_gen_1_s0_translator_avalon_anti_slave_0_writedata),  //           .writedata
		.avs_s0_readdata   (wave_gen_1_s0_translator_avalon_anti_slave_0_readdata),   //           .readdata
		.avs_s0_address    (wave_gen_1_s0_translator_avalon_anti_slave_0_address),    //           .address
		.clk_source        (nios_clk_clk),                                            // clk_source.clk
		.dac               (wave_gen_1_dac_export)                                    //        dac.export
	);

	wave_gen #(
		.AmpMax       (14'b11111111111111),
		.AmpMin       (14'b00000000000000),
		.FreqDiv      (34'b0000000000000000000000000000010100),
		.SamplePonint (13'b0000100000000)
	) wave_gen_2 (
		.clk               (altpll_0_c0_clk),                                         //      clock.clk
		.reset_n           (~rst_controller_001_reset_out_reset),                     //      reset.reset_n
		.avs_s0_chipselect (wave_gen_2_s0_translator_avalon_anti_slave_0_chipselect), //         s0.chipselect
		.avs_s0_write      (wave_gen_2_s0_translator_avalon_anti_slave_0_write),      //           .write
		.avs_s0_read       (wave_gen_2_s0_translator_avalon_anti_slave_0_read),       //           .read
		.avs_s0_writedata  (wave_gen_2_s0_translator_avalon_anti_slave_0_writedata),  //           .writedata
		.avs_s0_readdata   (wave_gen_2_s0_translator_avalon_anti_slave_0_readdata),   //           .readdata
		.avs_s0_address    (wave_gen_2_s0_translator_avalon_anti_slave_0_address),    //           .address
		.clk_source        (nios_clk_clk),                                            // clk_source.clk
		.dac               (wave_gen_2_dac_export)                                    //        dac.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (27),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (27),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_instruction_master_translator (
		.clk                      (nios_clk_clk),                                                                //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address              (nios2_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (nios2_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_byteenable            (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_write                 (1'b0),                                                                        //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.av_debugaccess           (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (27),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (27),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_data_master_translator (
		.clk                      (nios_clk_clk),                                                         //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address              (nios2_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios2_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2_data_master_read),                                               //                          .read
		.av_readdata              (nios2_data_master_readdata),                                           //                          .readdata
		.av_write                 (nios2_data_master_write),                                              //                          .write
		.av_writedata             (nios2_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                 //               (terminated)
		.av_begintransfer         (1'b0),                                                                 //               (terminated)
		.av_chipselect            (1'b0),                                                                 //               (terminated)
		.av_readdatavalid         (),                                                                     //               (terminated)
		.av_lock                  (1'b0),                                                                 //               (terminated)
		.uav_clken                (),                                                                     //               (terminated)
		.av_clken                 (1'b1),                                                                 //               (terminated)
		.uav_response             (2'b00),                                                                //               (terminated)
		.av_response              (),                                                                     //               (terminated)
		.uav_writeresponserequest (),                                                                     //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                 //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                 //               (terminated)
		.av_writeresponsevalid    ()                                                                      //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (27),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (27),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_0_read_master_translator (
		.clk                      (nios_clk_clk),                                                         //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address              (dma_0_read_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (dma_0_read_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (dma_0_read_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (dma_0_read_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (dma_0_read_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (dma_0_read_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (dma_0_read_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (dma_0_read_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (dma_0_read_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (dma_0_read_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (dma_0_read_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (dma_0_read_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (dma_0_read_master_waitrequest),                                        //                          .waitrequest
		.av_chipselect            (dma_0_read_master_chipselect),                                         //                          .chipselect
		.av_read                  (~dma_0_read_master_read),                                              //                          .read
		.av_readdata              (dma_0_read_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (dma_0_read_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                 //               (terminated)
		.av_byteenable            (4'b1111),                                                              //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                 //               (terminated)
		.av_begintransfer         (1'b0),                                                                 //               (terminated)
		.av_write                 (1'b0),                                                                 //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                 //               (terminated)
		.av_lock                  (1'b0),                                                                 //               (terminated)
		.av_debugaccess           (1'b0),                                                                 //               (terminated)
		.uav_clken                (),                                                                     //               (terminated)
		.av_clken                 (1'b1),                                                                 //               (terminated)
		.uav_response             (2'b00),                                                                //               (terminated)
		.av_response              (),                                                                     //               (terminated)
		.uav_writeresponserequest (),                                                                     //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                 //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                 //               (terminated)
		.av_writeresponsevalid    ()                                                                      //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_jtag_debug_module_translator (
		.clk                      (nios_clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address              (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                                   //              (terminated)
		.av_burstcount            (),                                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                                               //              (terminated)
		.av_writebyteenable       (),                                                                                   //              (terminated)
		.av_lock                  (),                                                                                   //              (terminated)
		.av_chipselect            (),                                                                                   //              (terminated)
		.av_clken                 (),                                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                                               //              (terminated)
		.av_outputenable          (),                                                                                   //              (terminated)
		.uav_response             (),                                                                                   //              (terminated)
		.av_response              (2'b00),                                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) epcs_flash_epcs_control_port_translator (
		.clk                      (nios_clk_clk),                                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                          //                    reset.reset
		.uav_address              (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                                        //              (terminated)
		.av_burstcount            (),                                                                                        //              (terminated)
		.av_byteenable            (),                                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                                        //              (terminated)
		.av_lock                  (),                                                                                        //              (terminated)
		.av_clken                 (),                                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                                    //              (terminated)
		.av_debugaccess           (),                                                                                        //              (terminated)
		.av_outputenable          (),                                                                                        //              (terminated)
		.uav_response             (),                                                                                        //              (terminated)
		.av_response              (2'b00),                                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_ram_s1_translator (
		.clk                      (nios_clk_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address              (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_ram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_ram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_ram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_ram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_ram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_ram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_ram_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (26),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_ddr2_clock_bridge_s0_translator (
		.clk                      (nios_clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address              (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (cpu_ddr2_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                                    //              (terminated)
		.av_lock                  (),                                                                                    //              (terminated)
		.av_chipselect            (),                                                                                    //              (terminated)
		.av_clken                 (),                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                //              (terminated)
		.av_outputenable          (),                                                                                    //              (terminated)
		.uav_response             (),                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) slow_peripheral_bridge_s0_translator (
		.clk                      (nios_clk_clk),                                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                       //                    reset.reset
		.uav_address              (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                     //              (terminated)
		.av_lock                  (),                                                                                     //              (terminated)
		.av_chipselect            (),                                                                                     //              (terminated)
		.av_clken                 (),                                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                                 //              (terminated)
		.av_outputenable          (),                                                                                     //              (terminated)
		.uav_response             (),                                                                                     //              (terminated)
		.av_response              (2'b00),                                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (27),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dma_0_control_port_slave_translator (
		.clk                      (nios_clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address              (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (dma_0_control_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (dma_0_control_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (dma_0_control_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (dma_0_control_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (dma_0_control_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                                    //              (terminated)
		.av_begintransfer         (),                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                    //              (terminated)
		.av_byteenable            (),                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                    //              (terminated)
		.av_lock                  (),                                                                                    //              (terminated)
		.av_clken                 (),                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                    //              (terminated)
		.uav_response             (),                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                 //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (10),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (10),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) slow_peripheral_bridge_m0_translator (
		.clk                      (altpll_0_c0_clk),                                                              //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                     reset.reset
		.uav_address              (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (slow_peripheral_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (slow_peripheral_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (slow_peripheral_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable            (slow_peripheral_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read                  (slow_peripheral_bridge_m0_read),                                               //                          .read
		.av_readdata              (slow_peripheral_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid         (slow_peripheral_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (slow_peripheral_bridge_m0_write),                                              //                          .write
		.av_writedata             (slow_peripheral_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess           (slow_peripheral_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer    (1'b0),                                                                         //               (terminated)
		.av_begintransfer         (1'b0),                                                                         //               (terminated)
		.av_chipselect            (1'b0),                                                                         //               (terminated)
		.av_lock                  (1'b0),                                                                         //               (terminated)
		.uav_clken                (),                                                                             //               (terminated)
		.av_clken                 (1'b1),                                                                         //               (terminated)
		.uav_response             (2'b00),                                                                        //               (terminated)
		.av_response              (),                                                                             //               (terminated)
		.uav_writeresponserequest (),                                                                             //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                         //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                         //               (terminated)
		.av_writeresponsevalid    ()                                                                              //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (10),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (10),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_0_write_master_translator (
		.clk                      (nios_clk_clk),                                                          //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                     reset.reset
		.uav_address              (dma_0_write_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (dma_0_write_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (dma_0_write_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (dma_0_write_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (dma_0_write_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (dma_0_write_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (dma_0_write_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (dma_0_write_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (dma_0_write_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (dma_0_write_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (dma_0_write_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (dma_0_write_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (dma_0_write_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (dma_0_write_master_byteenable),                                         //                          .byteenable
		.av_chipselect            (dma_0_write_master_chipselect),                                         //                          .chipselect
		.av_write                 (~dma_0_write_master_write),                                             //                          .write
		.av_writedata             (dma_0_write_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                  //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                  //               (terminated)
		.av_begintransfer         (1'b0),                                                                  //               (terminated)
		.av_read                  (1'b0),                                                                  //               (terminated)
		.av_readdata              (),                                                                      //               (terminated)
		.av_readdatavalid         (),                                                                      //               (terminated)
		.av_lock                  (1'b0),                                                                  //               (terminated)
		.av_debugaccess           (1'b0),                                                                  //               (terminated)
		.uav_clken                (),                                                                      //               (terminated)
		.av_clken                 (1'b1),                                                                  //               (terminated)
		.uav_response             (2'b00),                                                                 //               (terminated)
		.av_response              (),                                                                      //               (terminated)
		.uav_writeresponserequest (),                                                                      //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                  //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                  //               (terminated)
		.av_writeresponsevalid    ()                                                                       //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) altpll_0_pll_slave_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                            //                    reset.reset
		.uav_address              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (altpll_0_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (altpll_0_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (altpll_0_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_chipselect            (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                      (altpll_0_c0_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                             //                    reset.reset
		.uav_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                               //              (terminated)
		.av_read                  (),                                                                               //              (terminated)
		.av_writedata             (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                      (altpll_0_c0_clk),                                                                          //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                       //                    reset.reset
		.uav_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) systimer_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                        //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (systimer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (systimer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (systimer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (systimer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (systimer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (systimer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (systimer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (systimer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (systimer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (systimer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (systimer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (systimer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (systimer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (systimer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_key_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address              (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pio_key_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pio_key_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (pio_key_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pio_key_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pio_key_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) spi_0_spi_control_port_translator (
		.clk                      (altpll_0_c0_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                //                    reset.reset
		.uav_address              (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (spi_0_spi_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (spi_0_spi_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (spi_0_spi_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (spi_0_spi_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (spi_0_spi_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (spi_0_spi_control_port_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_byteenable            (),                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart_0_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                      //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                   //                    reset.reset
		.uav_address              (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (uart_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (uart_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (uart_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (uart_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (uart_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (uart_0_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect            (uart_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_led_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address              (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pio_led_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pio_led_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (pio_led_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pio_led_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pio_led_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timestamp_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timestamp_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timestamp_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timestamp_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timestamp_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timestamp_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) spi_ad5781_spi_control_port_translator (
		.clk                      (altpll_0_c0_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                     //                    reset.reset
		.uav_address              (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (spi_ad5781_spi_control_port_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ad9245_2_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                        //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read                  (ad9245_2_s1_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata              (ad9245_2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_chipselect            (ad9245_2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_address               (),                                                                       //              (terminated)
		.av_write                 (),                                                                       //              (terminated)
		.av_writedata             (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (5),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) clk_gen_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address              (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (clk_gen_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (clk_gen_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (clk_gen_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (clk_gen_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (clk_gen_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (clk_gen_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) oc_i2c_master_0_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                            //                    reset.reset
		.uav_address              (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_waitrequest           (~oc_i2c_master_0_s1_translator_avalon_anti_slave_0_waitrequest),                //                         .waitrequest
		.av_chipselect            (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) spi_master_0_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                         //                    reset.reset
		.uav_address              (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (spi_master_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (spi_master_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (spi_master_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (spi_master_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (spi_master_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (spi_master_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_burstcount            (),                                                                           //              (terminated)
		.av_byteenable            (),                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                       //              (terminated)
		.av_waitrequest           (1'b0),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_lock                  (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_debugaccess           (),                                                                           //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ad9266_spi_control_port_translator (
		.clk                      (altpll_0_c0_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ad9266_spi_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ad9266_spi_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ad9266_spi_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ad9266_spi_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ad9266_spi_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ad9266_spi_control_port_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                                   //              (terminated)
		.av_burstcount            (),                                                                                   //              (terminated)
		.av_byteenable            (),                                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                                               //              (terminated)
		.av_writebyteenable       (),                                                                                   //              (terminated)
		.av_lock                  (),                                                                                   //              (terminated)
		.av_clken                 (),                                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                                               //              (terminated)
		.av_debugaccess           (),                                                                                   //              (terminated)
		.av_outputenable          (),                                                                                   //              (terminated)
		.uav_response             (),                                                                                   //              (terminated)
		.av_response              (2'b00),                                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ad9245_1_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                        //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read                  (ad9245_1_s1_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata              (ad9245_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_chipselect            (ad9245_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_address               (),                                                                       //              (terminated)
		.av_write                 (),                                                                       //              (terminated)
		.av_writedata             (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dac2904_1_s0_translator (
		.clk                      (altpll_0_c0_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write                 (dac2904_1_s0_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata             (dac2904_1_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (dac2904_1_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (dac2904_1_s0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_address               (),                                                                        //              (terminated)
		.av_read                  (),                                                                        //              (terminated)
		.av_readdata              (32'b11011110101011011101111010101101),                                    //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dac2904_2_s0_translator (
		.clk                      (altpll_0_c0_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write                 (dac2904_2_s0_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata             (dac2904_2_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (dac2904_2_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (dac2904_2_s0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_address               (),                                                                        //              (terminated)
		.av_read                  (),                                                                        //              (terminated)
		.av_readdata              (32'b11011110101011011101111010101101),                                    //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dac2904_3_s0_translator (
		.clk                      (altpll_0_c0_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write                 (dac2904_3_s0_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata             (dac2904_3_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (dac2904_3_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (dac2904_3_s0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_address               (),                                                                        //              (terminated)
		.av_read                  (),                                                                        //              (terminated)
		.av_readdata              (32'b11011110101011011101111010101101),                                    //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dac2904_4_s0_translator (
		.clk                      (altpll_0_c0_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write                 (dac2904_4_s0_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata             (dac2904_4_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (dac2904_4_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (dac2904_4_s0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_address               (),                                                                        //              (terminated)
		.av_read                  (),                                                                        //              (terminated)
		.av_readdata              (32'b11011110101011011101111010101101),                                    //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) wave_gen_0_s0_translator (
		.clk                      (altpll_0_c0_clk),                                                          //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (wave_gen_0_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (wave_gen_0_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (wave_gen_0_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (wave_gen_0_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (wave_gen_0_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (wave_gen_0_s0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) demodulation_0_s0_translator (
		.clk                      (altpll_0_c0_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (demodulation_0_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (demodulation_0_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (demodulation_0_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (demodulation_0_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (demodulation_0_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (demodulation_0_s0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) wave_gen_1_s0_translator (
		.clk                      (altpll_0_c0_clk),                                                          //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (wave_gen_1_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (wave_gen_1_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (wave_gen_1_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (wave_gen_1_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (wave_gen_1_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (wave_gen_1_s0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) wave_gen_2_s0_translator (
		.clk                      (altpll_0_c0_clk),                                                          //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (wave_gen_2_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (wave_gen_2_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (wave_gen_2_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (wave_gen_2_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (wave_gen_2_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (wave_gen_2_s0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_ddr2_clock_bridge_m0_translator (
		.clk                      (ddr2_sysclk_clk),                                                             //                       clk.clk
		.reset                    (rst_controller_005_reset_out_reset),                                          //                     reset.reset
		.uav_address              (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_ddr2_clock_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_ddr2_clock_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (cpu_ddr2_clock_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable            (cpu_ddr2_clock_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read                  (cpu_ddr2_clock_bridge_m0_read),                                               //                          .read
		.av_readdata              (cpu_ddr2_clock_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid         (cpu_ddr2_clock_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (cpu_ddr2_clock_bridge_m0_write),                                              //                          .write
		.av_writedata             (cpu_ddr2_clock_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess           (cpu_ddr2_clock_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (24),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (3),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (5),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ddr2_s1_translator (
		.clk                      (ddr2_sysclk_clk),                                                    //                      clk.clk
		.reset                    (~ddr2_reset_request_n_reset),                                        //                    reset.reset
		.uav_address              (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ddr2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ddr2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ddr2_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ddr2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ddr2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_beginbursttransfer    (ddr2_s1_translator_avalon_anti_slave_0_beginbursttransfer),          //                         .beginbursttransfer
		.av_burstcount            (ddr2_s1_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (ddr2_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (ddr2_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (~ddr2_s1_translator_avalon_anti_slave_0_waitrequest),                //                         .waitrequest
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_chipselect            (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_BEGIN_BURST           (82),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.PKT_BURST_TYPE_H          (79),
		.PKT_BURST_TYPE_L          (78),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_TRANS_EXCLUSIVE       (68),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (87),
		.PKT_THREAD_ID_H           (90),
		.PKT_THREAD_ID_L           (90),
		.PKT_CACHE_H               (97),
		.PKT_CACHE_L               (94),
		.PKT_DATA_SIDEBAND_H       (81),
		.PKT_DATA_SIDEBAND_L       (81),
		.PKT_QOS_H                 (83),
		.PKT_QOS_L                 (83),
		.PKT_ADDR_SIDEBAND_H       (80),
		.PKT_ADDR_SIDEBAND_L       (80),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.ST_DATA_W                 (100),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (nios_clk_clk),                                                                         //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address              (nios2_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                                //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                                 //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                              //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                                        //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                          //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                                //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_BEGIN_BURST           (82),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.PKT_BURST_TYPE_H          (79),
		.PKT_BURST_TYPE_L          (78),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_TRANS_EXCLUSIVE       (68),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (87),
		.PKT_THREAD_ID_H           (90),
		.PKT_THREAD_ID_L           (90),
		.PKT_CACHE_H               (97),
		.PKT_CACHE_L               (94),
		.PKT_DATA_SIDEBAND_H       (81),
		.PKT_DATA_SIDEBAND_L       (81),
		.PKT_QOS_H                 (83),
		.PKT_QOS_L                 (83),
		.PKT_ADDR_SIDEBAND_H       (80),
		.PKT_ADDR_SIDEBAND_L       (80),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.ST_DATA_W                 (100),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (nios_clk_clk),                                                                  //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address              (nios2_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                    //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                     //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                  //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                              //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                    //          .ready
		.av_response             (),                                                                              // (terminated)
		.av_writeresponserequest (1'b0),                                                                          // (terminated)
		.av_writeresponsevalid   ()                                                                               // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_BEGIN_BURST           (82),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.PKT_BURST_TYPE_H          (79),
		.PKT_BURST_TYPE_L          (78),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_TRANS_EXCLUSIVE       (68),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (87),
		.PKT_THREAD_ID_H           (90),
		.PKT_THREAD_ID_L           (90),
		.PKT_CACHE_H               (97),
		.PKT_CACHE_L               (94),
		.PKT_DATA_SIDEBAND_H       (81),
		.PKT_DATA_SIDEBAND_L       (81),
		.PKT_QOS_H                 (83),
		.PKT_QOS_L                 (83),
		.PKT_ADDR_SIDEBAND_H       (80),
		.PKT_ADDR_SIDEBAND_L       (80),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.ST_DATA_W                 (100),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_0_read_master_translator_avalon_universal_master_0_agent (
		.clk                     (nios_clk_clk),                                                                  //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address              (dma_0_read_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (dma_0_read_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (dma_0_read_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (dma_0_read_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (dma_0_read_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (dma_0_read_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (dma_0_read_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (dma_0_read_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (dma_0_read_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (dma_0_read_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (dma_0_read_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_003_src2_valid),                                                 //        rp.valid
		.rp_data                 (rsp_xbar_demux_003_src2_data),                                                  //          .data
		.rp_channel              (rsp_xbar_demux_003_src2_channel),                                               //          .channel
		.rp_startofpacket        (rsp_xbar_demux_003_src2_startofpacket),                                         //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_003_src2_endofpacket),                                           //          .endofpacket
		.rp_ready                (rsp_xbar_demux_003_src2_ready),                                                 //          .ready
		.av_response             (),                                                                              // (terminated)
		.av_writeresponserequest (1'b0),                                                                          // (terminated)
		.av_writeresponsevalid   ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (100),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (nios_clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                     //                .channel
		.rf_sink_ready           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (101),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (nios_clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (100),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (nios_clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                    //       clk_reset.reset
		.m0_address              (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                                        //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                                        //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                         //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                                      //                .channel
		.rf_sink_ready           (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (101),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (nios_clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.in_data           (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (100),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_ram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (nios_clk_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                       //                .channel
		.rf_sink_ready           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (101),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (nios_clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (100),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (nios_clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                                  //                .channel
		.rf_sink_ready           (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (101),
		.FIFO_DEPTH          (73),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (nios_clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (100),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (nios_clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                                //                .channel
		.rf_sink_ready           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (101),
		.FIFO_DEPTH          (81),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (nios_clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (86),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (87),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (93),
		.PKT_PROTECTION_L          (91),
		.PKT_RESPONSE_STATUS_H     (99),
		.PKT_RESPONSE_STATUS_L     (98),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (100),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_0_control_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (nios_clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                               //                .channel
		.rf_sink_ready           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (101),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (nios_clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_BEGIN_BURST           (63),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.PKT_BURST_TYPE_H          (60),
		.PKT_BURST_TYPE_L          (59),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_TRANS_EXCLUSIVE       (51),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_THREAD_ID_H           (75),
		.PKT_THREAD_ID_L           (75),
		.PKT_CACHE_H               (82),
		.PKT_CACHE_L               (79),
		.PKT_DATA_SIDEBAND_H       (62),
		.PKT_DATA_SIDEBAND_L       (62),
		.PKT_QOS_H                 (64),
		.PKT_QOS_L                 (64),
		.PKT_ADDR_SIDEBAND_H       (61),
		.PKT_ADDR_SIDEBAND_L       (61),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.ST_DATA_W                 (85),
		.ST_CHANNEL_W              (24),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                       //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.av_address              (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_001_rsp_src_valid),                                                             //        rp.valid
		.rp_data                 (limiter_001_rsp_src_data),                                                              //          .data
		.rp_channel              (limiter_001_rsp_src_channel),                                                           //          .channel
		.rp_startofpacket        (limiter_001_rsp_src_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket          (limiter_001_rsp_src_endofpacket),                                                       //          .endofpacket
		.rp_ready                (limiter_001_rsp_src_ready),                                                             //          .ready
		.av_response             (),                                                                                      // (terminated)
		.av_writeresponserequest (1'b0),                                                                                  // (terminated)
		.av_writeresponsevalid   ()                                                                                       // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_BEGIN_BURST           (63),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.PKT_BURST_TYPE_H          (60),
		.PKT_BURST_TYPE_L          (59),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_TRANS_EXCLUSIVE       (51),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_THREAD_ID_H           (75),
		.PKT_THREAD_ID_L           (75),
		.PKT_CACHE_H               (82),
		.PKT_CACHE_L               (79),
		.PKT_DATA_SIDEBAND_H       (62),
		.PKT_DATA_SIDEBAND_L       (62),
		.PKT_QOS_H                 (64),
		.PKT_QOS_L                 (64),
		.PKT_ADDR_SIDEBAND_H       (61),
		.PKT_ADDR_SIDEBAND_L       (61),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.ST_DATA_W                 (85),
		.ST_CHANNEL_W              (24),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_0_write_master_translator_avalon_universal_master_0_agent (
		.clk                     (nios_clk_clk),                                                                   //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.av_address              (dma_0_write_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (dma_0_write_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (dma_0_write_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (dma_0_write_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (dma_0_write_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (dma_0_write_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (dma_0_write_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (dma_0_write_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (dma_0_write_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (dma_0_write_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (dma_0_write_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_004_src_valid),                                                     //        rp.valid
		.rp_data                 (rsp_xbar_mux_004_src_data),                                                      //          .data
		.rp_channel              (rsp_xbar_mux_004_src_channel),                                                   //          .channel
		.rp_startofpacket        (rsp_xbar_mux_004_src_startofpacket),                                             //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_004_src_endofpacket),                                               //          .endofpacket
		.rp_ready                (rsp_xbar_mux_004_src_ready),                                                     //          .ready
		.av_response             (),                                                                               // (terminated)
		.av_writeresponserequest (1'b0),                                                                           // (terminated)
		.av_writeresponsevalid   ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                       //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                       //                .valid
		.cp_data                 (crosser_out_data),                                                                        //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                     //                .channel
		.rf_sink_ready           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                // clk_reset.reset
		.in_data           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_startofpacket  (1'b0),                                                                              // (terminated)
		.in_endofpacket    (1'b0),                                                                              // (terminated)
		.out_startofpacket (),                                                                                  // (terminated)
		.out_endofpacket   (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src1_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src1_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_003_src1_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src1_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src1_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src1_channel),                                                          //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_startofpacket  (1'b0),                                                                               // (terminated)
		.in_endofpacket    (1'b0),                                                                               // (terminated)
		.out_startofpacket (),                                                                                   // (terminated)
		.out_endofpacket   (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src2_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src2_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_003_src2_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src2_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src2_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src2_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                                         // (terminated)
		.out_startofpacket (),                                                                                             // (terminated)
		.out_endofpacket   (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) systimer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (systimer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (systimer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (systimer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (systimer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (systimer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (systimer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (systimer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (systimer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (systimer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (systimer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (systimer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (systimer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (systimer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (systimer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src3_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src3_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_003_src3_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src3_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src3_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src3_channel),                                                  //                .channel
		.rf_sink_ready           (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.in_data           (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                       // (terminated)
		.out_startofpacket (),                                                                           // (terminated)
		.out_endofpacket   (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pio_key_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src4_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src4_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_003_src4_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src4_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src4_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src4_channel),                                                 //                .channel
		.rf_sink_ready           (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.in_data           (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                     // (terminated)
		.csr_read          (1'b0),                                                                      // (terminated)
		.csr_write         (1'b0),                                                                      // (terminated)
		.csr_readdata      (),                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                      // (terminated)
		.almost_full_data  (),                                                                          // (terminated)
		.almost_empty_data (),                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                      // (terminated)
		.out_startofpacket (),                                                                          // (terminated)
		.out_endofpacket   (),                                                                          // (terminated)
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_channel        (1'b0),                                                                      // (terminated)
		.out_channel       ()                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) spi_0_spi_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src5_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src5_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_003_src5_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src5_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src5_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src5_channel),                                                             //                .channel
		.rf_sink_ready           (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_startofpacket  (1'b0),                                                                                  // (terminated)
		.in_endofpacket    (1'b0),                                                                                  // (terminated)
		.out_startofpacket (),                                                                                      // (terminated)
		.out_endofpacket   (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) uart_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src6_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src6_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_003_src6_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src6_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src6_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src6_channel),                                                //                .channel
		.rf_sink_ready           (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.in_data           (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                    // (terminated)
		.csr_read          (1'b0),                                                                     // (terminated)
		.csr_write         (1'b0),                                                                     // (terminated)
		.csr_readdata      (),                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                     // (terminated)
		.almost_full_data  (),                                                                         // (terminated)
		.almost_empty_data (),                                                                         // (terminated)
		.in_startofpacket  (1'b0),                                                                     // (terminated)
		.in_endofpacket    (1'b0),                                                                     // (terminated)
		.out_startofpacket (),                                                                         // (terminated)
		.out_endofpacket   (),                                                                         // (terminated)
		.in_empty          (1'b0),                                                                     // (terminated)
		.out_empty         (),                                                                         // (terminated)
		.in_error          (1'b0),                                                                     // (terminated)
		.out_error         (),                                                                         // (terminated)
		.in_channel        (1'b0),                                                                     // (terminated)
		.out_channel       ()                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pio_led_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src7_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src7_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_003_src7_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src7_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src7_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src7_channel),                                                 //                .channel
		.rf_sink_ready           (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.in_data           (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                     // (terminated)
		.csr_read          (1'b0),                                                                      // (terminated)
		.csr_write         (1'b0),                                                                      // (terminated)
		.csr_readdata      (),                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                      // (terminated)
		.almost_full_data  (),                                                                          // (terminated)
		.almost_empty_data (),                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                      // (terminated)
		.out_startofpacket (),                                                                          // (terminated)
		.out_endofpacket   (),                                                                          // (terminated)
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_channel        (1'b0),                                                                      // (terminated)
		.out_channel       ()                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timestamp_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src8_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src8_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_003_src8_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src8_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src8_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src8_channel),                                                   //                .channel
		.rf_sink_ready           (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_startofpacket  (1'b0),                                                                        // (terminated)
		.in_endofpacket    (1'b0),                                                                        // (terminated)
		.out_startofpacket (),                                                                            // (terminated)
		.out_endofpacket   (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src9_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src9_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_003_src9_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src9_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src9_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src9_channel),                                                                  //                .channel
		.rf_sink_ready           (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                                       // (terminated)
		.out_startofpacket (),                                                                                           // (terminated)
		.out_endofpacket   (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ad9245_2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ad9245_2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src10_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src10_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_003_src10_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src10_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src10_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src10_channel),                                                 //                .channel
		.rf_sink_ready           (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.in_data           (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                       // (terminated)
		.out_startofpacket (),                                                                           // (terminated)
		.out_endofpacket   (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) clk_gen_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (clk_gen_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (clk_gen_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (clk_gen_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (clk_gen_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (clk_gen_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (clk_gen_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src11_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src11_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_003_src11_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src11_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src11_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src11_channel),                                                //                .channel
		.rf_sink_ready           (clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (clk_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (clk_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (clk_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (clk_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (clk_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (clk_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (clk_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (clk_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (clk_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (clk_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (clk_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.in_data           (clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (clk_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                     // (terminated)
		.csr_read          (1'b0),                                                                      // (terminated)
		.csr_write         (1'b0),                                                                      // (terminated)
		.csr_readdata      (),                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                      // (terminated)
		.almost_full_data  (),                                                                          // (terminated)
		.almost_empty_data (),                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                      // (terminated)
		.out_startofpacket (),                                                                          // (terminated)
		.out_endofpacket   (),                                                                          // (terminated)
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_channel        (1'b0),                                                                      // (terminated)
		.out_channel       ()                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src12_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src12_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_003_src12_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src12_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src12_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src12_channel),                                                        //                .channel
		.rf_sink_ready           (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_startofpacket  (1'b0),                                                                              // (terminated)
		.in_endofpacket    (1'b0),                                                                              // (terminated)
		.out_startofpacket (),                                                                                  // (terminated)
		.out_endofpacket   (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) spi_master_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (spi_master_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src13_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src13_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_003_src13_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src13_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src13_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src13_channel),                                                     //                .channel
		.rf_sink_ready           (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_startofpacket  (1'b0),                                                                           // (terminated)
		.in_endofpacket    (1'b0),                                                                           // (terminated)
		.out_startofpacket (),                                                                               // (terminated)
		.out_endofpacket   (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ad9266_spi_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src14_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src14_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_003_src14_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src14_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src14_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src14_channel),                                                             //                .channel
		.rf_sink_ready           (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_startofpacket  (1'b0),                                                                                   // (terminated)
		.in_endofpacket    (1'b0),                                                                                   // (terminated)
		.out_startofpacket (),                                                                                       // (terminated)
		.out_endofpacket   (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ad9245_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ad9245_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_021_src_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_021_src_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_021_src_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_021_src_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_021_src_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_021_src_channel),                                                     //                .channel
		.rf_sink_ready           (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.in_data           (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                       // (terminated)
		.out_startofpacket (),                                                                           // (terminated)
		.out_endofpacket   (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dac2904_1_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dac2904_1_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_022_src_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_mux_022_src_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_mux_022_src_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_mux_022_src_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_022_src_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_mux_022_src_channel),                                                      //                .channel
		.rf_sink_ready           (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_startofpacket  (1'b0),                                                                        // (terminated)
		.in_endofpacket    (1'b0),                                                                        // (terminated)
		.out_startofpacket (),                                                                            // (terminated)
		.out_endofpacket   (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dac2904_2_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dac2904_2_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src17_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src17_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_003_src17_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src17_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src17_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src17_channel),                                                  //                .channel
		.rf_sink_ready           (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_startofpacket  (1'b0),                                                                        // (terminated)
		.in_endofpacket    (1'b0),                                                                        // (terminated)
		.out_startofpacket (),                                                                            // (terminated)
		.out_endofpacket   (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dac2904_3_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dac2904_3_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src18_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src18_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_003_src18_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src18_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src18_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src18_channel),                                                  //                .channel
		.rf_sink_ready           (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_startofpacket  (1'b0),                                                                        // (terminated)
		.in_endofpacket    (1'b0),                                                                        // (terminated)
		.out_startofpacket (),                                                                            // (terminated)
		.out_endofpacket   (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dac2904_4_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dac2904_4_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src19_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src19_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_003_src19_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src19_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src19_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src19_channel),                                                  //                .channel
		.rf_sink_ready           (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_startofpacket  (1'b0),                                                                        // (terminated)
		.in_endofpacket    (1'b0),                                                                        // (terminated)
		.out_startofpacket (),                                                                            // (terminated)
		.out_endofpacket   (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) wave_gen_0_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src20_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src20_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_003_src20_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src20_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src20_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src20_channel),                                                   //                .channel
		.rf_sink_ready           (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                         // (terminated)
		.out_startofpacket (),                                                                             // (terminated)
		.out_endofpacket   (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) demodulation_0_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (demodulation_0_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src21_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src21_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_003_src21_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src21_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src21_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src21_channel),                                                       //                .channel
		.rf_sink_ready           (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_startofpacket  (1'b0),                                                                             // (terminated)
		.in_endofpacket    (1'b0),                                                                             // (terminated)
		.out_startofpacket (),                                                                                 // (terminated)
		.out_endofpacket   (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) wave_gen_1_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src22_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src22_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_003_src22_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src22_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src22_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src22_channel),                                                   //                .channel
		.rf_sink_ready           (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                         // (terminated)
		.out_startofpacket (),                                                                             // (terminated)
		.out_endofpacket   (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (24),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) wave_gen_2_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src23_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src23_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_003_src23_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src23_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src23_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src23_channel),                                                   //                .channel
		.rf_sink_ready           (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                         // (terminated)
		.out_startofpacket (),                                                                             // (terminated)
		.out_endofpacket   (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.PKT_BURST_TYPE_H          (78),
		.PKT_BURST_TYPE_L          (77),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (84),
		.PKT_THREAD_ID_H           (85),
		.PKT_THREAD_ID_L           (85),
		.PKT_CACHE_H               (92),
		.PKT_CACHE_L               (89),
		.PKT_DATA_SIDEBAND_H       (80),
		.PKT_DATA_SIDEBAND_L       (80),
		.PKT_QOS_H                 (82),
		.PKT_QOS_L                 (82),
		.PKT_ADDR_SIDEBAND_H       (79),
		.PKT_ADDR_SIDEBAND_L       (79),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.ST_DATA_W                 (95),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk                     (ddr2_sysclk_clk),                                                                      //       clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                                   // clk_reset.reset
		.av_address              (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_030_src0_valid),                                                        //        rp.valid
		.rp_data                 (rsp_xbar_demux_030_src0_data),                                                         //          .data
		.rp_channel              (rsp_xbar_demux_030_src0_channel),                                                      //          .channel
		.rp_startofpacket        (rsp_xbar_demux_030_src0_startofpacket),                                                //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_030_src0_endofpacket),                                                  //          .endofpacket
		.rp_ready                (rsp_xbar_demux_030_src0_ready),                                                        //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (83),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (84),
		.PKT_DEST_ID_L             (84),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (73),
		.PKT_BYTE_CNT_H            (72),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (88),
		.PKT_PROTECTION_L          (86),
		.PKT_RESPONSE_STATUS_H     (94),
		.PKT_RESPONSE_STATUS_L     (93),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (95),
		.AVS_BURSTCOUNT_W          (5),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ddr2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (ddr2_sysclk_clk),                                                              //             clk.clk
		.reset                   (~ddr2_reset_request_n_reset),                                                  //       clk_reset.reset
		.m0_address              (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ddr2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ddr2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ddr2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ddr2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ddr2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ddr2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_005_src0_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_005_src0_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_005_src0_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_005_src0_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_005_src0_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_005_src0_channel),                                              //                .channel
		.rf_sink_ready           (ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ddr2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ddr2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ddr2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ddr2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ddr2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ddr2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ddr2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ddr2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ddr2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ddr2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ddr2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (96),
		.FIFO_DEPTH          (33),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (ddr2_sysclk_clk),                                                              //       clk.clk
		.reset             (~ddr2_reset_request_n_reset),                                                  // clk_reset.reset
		.in_data           (ddr2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ddr2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ddr2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ddr2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ddr2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ddr2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	nios2_addr_router addr_router (
		.sink_ready         (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (nios_clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_src_valid),                                                                //          .valid
		.src_data           (addr_router_src_data),                                                                 //          .data
		.src_channel        (addr_router_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                           //          .endofpacket
	);

	nios2_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (nios_clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                     //          .valid
		.src_data           (addr_router_001_src_data),                                                      //          .data
		.src_channel        (addr_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                //          .endofpacket
	);

	nios2_addr_router_002 addr_router_002 (
		.sink_ready         (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (nios_clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                     //          .valid
		.src_data           (addr_router_002_src_data),                                                      //          .data
		.src_channel        (addr_router_002_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                //          .endofpacket
	);

	nios2_id_router id_router (
		.sink_ready         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (nios_clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                //       src.ready
		.src_valid          (id_router_src_valid),                                                                //          .valid
		.src_data           (id_router_src_data),                                                                 //          .data
		.src_channel        (id_router_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                           //          .endofpacket
	);

	nios2_id_router id_router_001 (
		.sink_ready         (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (nios_clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                                 //       src.ready
		.src_valid          (id_router_001_src_valid),                                                                 //          .valid
		.src_data           (id_router_001_src_data),                                                                  //          .data
		.src_channel        (id_router_001_src_channel),                                                               //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                            //          .endofpacket
	);

	nios2_id_router id_router_002 (
		.sink_ready         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (nios_clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                  //       src.ready
		.src_valid          (id_router_002_src_valid),                                                  //          .valid
		.src_data           (id_router_002_src_data),                                                   //          .data
		.src_channel        (id_router_002_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                             //          .endofpacket
	);

	nios2_id_router_003 id_router_003 (
		.sink_ready         (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_ddr2_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (nios_clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                             //       src.ready
		.src_valid          (id_router_003_src_valid),                                                             //          .valid
		.src_data           (id_router_003_src_data),                                                              //          .data
		.src_channel        (id_router_003_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                        //          .endofpacket
	);

	nios2_id_router_004 id_router_004 (
		.sink_ready         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (nios_clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                              //       src.ready
		.src_valid          (id_router_004_src_valid),                                                              //          .valid
		.src_data           (id_router_004_src_data),                                                               //          .data
		.src_channel        (id_router_004_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                         //          .endofpacket
	);

	nios2_id_router_004 id_router_005 (
		.sink_ready         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (nios_clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                             //       src.ready
		.src_valid          (id_router_005_src_valid),                                                             //          .valid
		.src_data           (id_router_005_src_data),                                                              //          .data
		.src_channel        (id_router_005_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                        //          .endofpacket
	);

	nios2_addr_router_003 addr_router_003 (
		.sink_ready         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                             //          .valid
		.src_data           (addr_router_003_src_data),                                                              //          .data
		.src_channel        (addr_router_003_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                        //          .endofpacket
	);

	nios2_addr_router_004 addr_router_004 (
		.sink_ready         (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (nios_clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                      //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                      //          .valid
		.src_data           (addr_router_004_src_data),                                                       //          .data
		.src_channel        (addr_router_004_src_channel),                                                    //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                 //          .endofpacket
	);

	nios2_id_router_006 id_router_006 (
		.sink_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                       //       src.ready
		.src_valid          (id_router_006_src_valid),                                                       //          .valid
		.src_data           (id_router_006_src_data),                                                        //          .data
		.src_channel        (id_router_006_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                  //          .endofpacket
	);

	nios2_id_router_006 id_router_007 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                        //       src.ready
		.src_valid          (id_router_007_src_valid),                                                        //          .valid
		.src_data           (id_router_007_src_data),                                                         //          .data
		.src_channel        (id_router_007_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                   //          .endofpacket
	);

	nios2_id_router_006 id_router_008 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                  //          .valid
		.src_data           (id_router_008_src_data),                                                                   //          .data
		.src_channel        (id_router_008_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                             //          .endofpacket
	);

	nios2_id_router_006 id_router_009 (
		.sink_ready         (systimer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (systimer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (systimer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (systimer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (systimer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                //       src.ready
		.src_valid          (id_router_009_src_valid),                                                //          .valid
		.src_data           (id_router_009_src_data),                                                 //          .data
		.src_channel        (id_router_009_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                           //          .endofpacket
	);

	nios2_id_router_006 id_router_010 (
		.sink_ready         (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                               //       src.ready
		.src_valid          (id_router_010_src_valid),                                               //          .valid
		.src_data           (id_router_010_src_data),                                                //          .data
		.src_channel        (id_router_010_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                          //          .endofpacket
	);

	nios2_id_router_006 id_router_011 (
		.sink_ready         (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (spi_0_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                           //       src.ready
		.src_valid          (id_router_011_src_valid),                                                           //          .valid
		.src_data           (id_router_011_src_data),                                                            //          .data
		.src_channel        (id_router_011_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                      //          .endofpacket
	);

	nios2_id_router_006 id_router_012 (
		.sink_ready         (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                              //       src.ready
		.src_valid          (id_router_012_src_valid),                                              //          .valid
		.src_data           (id_router_012_src_data),                                               //          .data
		.src_channel        (id_router_012_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                         //          .endofpacket
	);

	nios2_id_router_006 id_router_013 (
		.sink_ready         (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                               //       src.ready
		.src_valid          (id_router_013_src_valid),                                               //          .valid
		.src_data           (id_router_013_src_data),                                                //          .data
		.src_channel        (id_router_013_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                          //          .endofpacket
	);

	nios2_id_router_006 id_router_014 (
		.sink_ready         (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                 //       src.ready
		.src_valid          (id_router_014_src_valid),                                                 //          .valid
		.src_data           (id_router_014_src_data),                                                  //          .data
		.src_channel        (id_router_014_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                            //          .endofpacket
	);

	nios2_id_router_006 id_router_015 (
		.sink_ready         (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (spi_ad5781_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                                //       src.ready
		.src_valid          (id_router_015_src_valid),                                                                //          .valid
		.src_data           (id_router_015_src_data),                                                                 //          .data
		.src_channel        (id_router_015_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                                           //          .endofpacket
	);

	nios2_id_router_006 id_router_016 (
		.sink_ready         (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ad9245_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                //       src.ready
		.src_valid          (id_router_016_src_valid),                                                //          .valid
		.src_data           (id_router_016_src_data),                                                 //          .data
		.src_channel        (id_router_016_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                           //          .endofpacket
	);

	nios2_id_router_006 id_router_017 (
		.sink_ready         (clk_gen_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (clk_gen_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (clk_gen_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (clk_gen_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (clk_gen_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                               //       src.ready
		.src_valid          (id_router_017_src_valid),                                               //          .valid
		.src_data           (id_router_017_src_data),                                                //          .data
		.src_channel        (id_router_017_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                          //          .endofpacket
	);

	nios2_id_router_006 id_router_018 (
		.sink_ready         (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                       //       src.ready
		.src_valid          (id_router_018_src_valid),                                                       //          .valid
		.src_data           (id_router_018_src_data),                                                        //          .data
		.src_channel        (id_router_018_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                                  //          .endofpacket
	);

	nios2_id_router_006 id_router_019 (
		.sink_ready         (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (spi_master_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                                    //       src.ready
		.src_valid          (id_router_019_src_valid),                                                    //          .valid
		.src_data           (id_router_019_src_data),                                                     //          .data
		.src_channel        (id_router_019_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                               //          .endofpacket
	);

	nios2_id_router_006 id_router_020 (
		.sink_ready         (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ad9266_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                                            //       src.ready
		.src_valid          (id_router_020_src_valid),                                                            //          .valid
		.src_data           (id_router_020_src_data),                                                             //          .data
		.src_channel        (id_router_020_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                                       //          .endofpacket
	);

	nios2_id_router_021 id_router_021 (
		.sink_ready         (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ad9245_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                                //       src.ready
		.src_valid          (id_router_021_src_valid),                                                //          .valid
		.src_data           (id_router_021_src_data),                                                 //          .data
		.src_channel        (id_router_021_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                           //          .endofpacket
	);

	nios2_id_router_021 id_router_022 (
		.sink_ready         (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dac2904_1_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                                                 //       src.ready
		.src_valid          (id_router_022_src_valid),                                                 //          .valid
		.src_data           (id_router_022_src_data),                                                  //          .data
		.src_channel        (id_router_022_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)                                            //          .endofpacket
	);

	nios2_id_router_006 id_router_023 (
		.sink_ready         (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dac2904_2_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_023_src_ready),                                                 //       src.ready
		.src_valid          (id_router_023_src_valid),                                                 //          .valid
		.src_data           (id_router_023_src_data),                                                  //          .data
		.src_channel        (id_router_023_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_023_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_023_src_endofpacket)                                            //          .endofpacket
	);

	nios2_id_router_006 id_router_024 (
		.sink_ready         (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dac2904_3_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_024_src_ready),                                                 //       src.ready
		.src_valid          (id_router_024_src_valid),                                                 //          .valid
		.src_data           (id_router_024_src_data),                                                  //          .data
		.src_channel        (id_router_024_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_024_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_024_src_endofpacket)                                            //          .endofpacket
	);

	nios2_id_router_006 id_router_025 (
		.sink_ready         (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dac2904_4_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_025_src_ready),                                                 //       src.ready
		.src_valid          (id_router_025_src_valid),                                                 //          .valid
		.src_data           (id_router_025_src_data),                                                  //          .data
		.src_channel        (id_router_025_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_025_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_025_src_endofpacket)                                            //          .endofpacket
	);

	nios2_id_router_006 id_router_026 (
		.sink_ready         (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (wave_gen_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_026_src_ready),                                                  //       src.ready
		.src_valid          (id_router_026_src_valid),                                                  //          .valid
		.src_data           (id_router_026_src_data),                                                   //          .data
		.src_channel        (id_router_026_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_026_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_026_src_endofpacket)                                             //          .endofpacket
	);

	nios2_id_router_006 id_router_027 (
		.sink_ready         (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (demodulation_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_027_src_ready),                                                      //       src.ready
		.src_valid          (id_router_027_src_valid),                                                      //          .valid
		.src_data           (id_router_027_src_data),                                                       //          .data
		.src_channel        (id_router_027_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_027_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_027_src_endofpacket)                                                 //          .endofpacket
	);

	nios2_id_router_006 id_router_028 (
		.sink_ready         (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (wave_gen_1_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_028_src_ready),                                                  //       src.ready
		.src_valid          (id_router_028_src_valid),                                                  //          .valid
		.src_data           (id_router_028_src_data),                                                   //          .data
		.src_channel        (id_router_028_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_028_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_028_src_endofpacket)                                             //          .endofpacket
	);

	nios2_id_router_006 id_router_029 (
		.sink_ready         (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (wave_gen_2_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_029_src_ready),                                                  //       src.ready
		.src_valid          (id_router_029_src_valid),                                                  //          .valid
		.src_data           (id_router_029_src_data),                                                   //          .data
		.src_channel        (id_router_029_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_029_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_029_src_endofpacket)                                             //          .endofpacket
	);

	nios2_addr_router_005 addr_router_005 (
		.sink_ready         (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_ddr2_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ddr2_sysclk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                            //          .valid
		.src_data           (addr_router_005_src_data),                                                             //          .data
		.src_channel        (addr_router_005_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                                       //          .endofpacket
	);

	nios2_id_router_030 id_router_030 (
		.sink_ready         (ddr2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ddr2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ddr2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ddr2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ddr2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (ddr2_sysclk_clk),                                                    //       clk.clk
		.reset              (~ddr2_reset_request_n_reset),                                        // clk_reset.reset
		.src_ready          (id_router_030_src_ready),                                            //       src.ready
		.src_valid          (id_router_030_src_valid),                                            //          .valid
		.src_data           (id_router_030_src_data),                                             //          .data
		.src_channel        (id_router_030_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_030_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_030_src_endofpacket)                                       //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (89),
		.PKT_DEST_ID_L             (87),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.MAX_OUTSTANDING_RESPONSES (72),
		.PIPELINED                 (0),
		.ST_DATA_W                 (100),
		.ST_CHANNEL_W              (6),
		.VALID_WIDTH               (6),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (nios_clk_clk),                   //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.MAX_OUTSTANDING_RESPONSES (5),
		.PIPELINED                 (0),
		.ST_DATA_W                 (85),
		.ST_CHANNEL_W              (24),
		.VALID_WIDTH               (24),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (altpll_0_c0_clk),                    //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_003_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_003_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_003_src_data),           //          .data
		.cmd_sink_channel       (addr_router_003_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_003_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_003_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_003_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_003_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_003_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_003_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_003_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_003_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (~ddr2_reset_request_n_reset),         // reset_in2.reset
		.clk        (nios_clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (~ddr2_reset_request_n_reset),         // reset_in2.reset
		.clk        (altpll_0_c0_clk),                     //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (~ddr2_reset_request_n_reset),         // reset_in2.reset
		.clk        (altpll_0_c1_clk),                     //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_003 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (altpll_0_c1_clk),                    //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_004 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (~ddr2_reset_request_n_reset),         // reset_in2.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_004_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (3),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_005 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2  (~ddr2_reset_request_n_reset),         // reset_in2.reset
		.clk        (ddr2_sysclk_clk),                     //       clk.clk
		.reset_out  (rst_controller_005_reset_out_reset),  // reset_out.reset
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	nios2_cmd_xbar_demux cmd_xbar_demux (
		.clk                (nios_clk_clk),                      //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket)    //           .endofpacket
	);

	nios2_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (nios_clk_clk),                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //          .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //      src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (nios_clk_clk),                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (nios_clk_clk),                          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (nios_clk_clk),                          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (nios_clk_clk),                          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_mux_003 cmd_xbar_mux_003 (
		.clk                 (nios_clk_clk),                          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux rsp_xbar_demux (
		.clk                (nios_clk_clk),                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (nios_clk_clk),                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (nios_clk_clk),                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (nios_clk_clk),                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_003_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_003_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_003_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_003_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_003_src2_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (nios_clk_clk),                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_demux_002 rsp_xbar_demux_005 (
		.clk                (nios_clk_clk),                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (nios_clk_clk),                          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (nios_clk_clk),                          //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_demux_003 cmd_xbar_demux_003 (
		.clk                 (altpll_0_c0_clk),                        //        clk.clk
		.reset               (rst_controller_001_reset_out_reset),     //  clk_reset.reset
		.sink_ready          (limiter_001_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_001_cmd_src_channel),            //           .channel
		.sink_data           (limiter_001_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_001_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_001_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_001_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_003_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_003_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_003_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_003_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_003_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_003_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_003_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_003_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_003_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_003_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_003_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_003_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_003_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_003_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_003_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_003_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_003_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_003_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_003_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_003_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_003_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_003_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_003_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_003_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_003_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_003_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_003_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_003_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_003_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_003_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_003_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_003_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_003_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_003_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_003_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_003_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_003_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_003_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_003_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_003_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_003_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_003_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_003_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_003_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_003_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_003_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_003_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_003_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_003_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_003_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_003_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_003_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_003_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_003_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_003_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_003_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_003_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_003_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_003_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_003_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_003_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_003_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_003_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_003_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_003_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_003_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_003_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_003_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_003_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_003_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_003_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_003_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_003_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_003_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_003_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_003_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_003_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_003_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_003_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_003_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_003_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_003_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_003_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_003_src13_endofpacket),   //           .endofpacket
		.src14_ready         (cmd_xbar_demux_003_src14_ready),         //      src14.ready
		.src14_valid         (cmd_xbar_demux_003_src14_valid),         //           .valid
		.src14_data          (cmd_xbar_demux_003_src14_data),          //           .data
		.src14_channel       (cmd_xbar_demux_003_src14_channel),       //           .channel
		.src14_startofpacket (cmd_xbar_demux_003_src14_startofpacket), //           .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_003_src14_endofpacket),   //           .endofpacket
		.src15_ready         (cmd_xbar_demux_003_src15_ready),         //      src15.ready
		.src15_valid         (cmd_xbar_demux_003_src15_valid),         //           .valid
		.src15_data          (cmd_xbar_demux_003_src15_data),          //           .data
		.src15_channel       (cmd_xbar_demux_003_src15_channel),       //           .channel
		.src15_startofpacket (cmd_xbar_demux_003_src15_startofpacket), //           .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_003_src15_endofpacket),   //           .endofpacket
		.src16_ready         (cmd_xbar_demux_003_src16_ready),         //      src16.ready
		.src16_valid         (cmd_xbar_demux_003_src16_valid),         //           .valid
		.src16_data          (cmd_xbar_demux_003_src16_data),          //           .data
		.src16_channel       (cmd_xbar_demux_003_src16_channel),       //           .channel
		.src16_startofpacket (cmd_xbar_demux_003_src16_startofpacket), //           .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_003_src16_endofpacket),   //           .endofpacket
		.src17_ready         (cmd_xbar_demux_003_src17_ready),         //      src17.ready
		.src17_valid         (cmd_xbar_demux_003_src17_valid),         //           .valid
		.src17_data          (cmd_xbar_demux_003_src17_data),          //           .data
		.src17_channel       (cmd_xbar_demux_003_src17_channel),       //           .channel
		.src17_startofpacket (cmd_xbar_demux_003_src17_startofpacket), //           .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_003_src17_endofpacket),   //           .endofpacket
		.src18_ready         (cmd_xbar_demux_003_src18_ready),         //      src18.ready
		.src18_valid         (cmd_xbar_demux_003_src18_valid),         //           .valid
		.src18_data          (cmd_xbar_demux_003_src18_data),          //           .data
		.src18_channel       (cmd_xbar_demux_003_src18_channel),       //           .channel
		.src18_startofpacket (cmd_xbar_demux_003_src18_startofpacket), //           .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_003_src18_endofpacket),   //           .endofpacket
		.src19_ready         (cmd_xbar_demux_003_src19_ready),         //      src19.ready
		.src19_valid         (cmd_xbar_demux_003_src19_valid),         //           .valid
		.src19_data          (cmd_xbar_demux_003_src19_data),          //           .data
		.src19_channel       (cmd_xbar_demux_003_src19_channel),       //           .channel
		.src19_startofpacket (cmd_xbar_demux_003_src19_startofpacket), //           .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_003_src19_endofpacket),   //           .endofpacket
		.src20_ready         (cmd_xbar_demux_003_src20_ready),         //      src20.ready
		.src20_valid         (cmd_xbar_demux_003_src20_valid),         //           .valid
		.src20_data          (cmd_xbar_demux_003_src20_data),          //           .data
		.src20_channel       (cmd_xbar_demux_003_src20_channel),       //           .channel
		.src20_startofpacket (cmd_xbar_demux_003_src20_startofpacket), //           .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_003_src20_endofpacket),   //           .endofpacket
		.src21_ready         (cmd_xbar_demux_003_src21_ready),         //      src21.ready
		.src21_valid         (cmd_xbar_demux_003_src21_valid),         //           .valid
		.src21_data          (cmd_xbar_demux_003_src21_data),          //           .data
		.src21_channel       (cmd_xbar_demux_003_src21_channel),       //           .channel
		.src21_startofpacket (cmd_xbar_demux_003_src21_startofpacket), //           .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_003_src21_endofpacket),   //           .endofpacket
		.src22_ready         (cmd_xbar_demux_003_src22_ready),         //      src22.ready
		.src22_valid         (cmd_xbar_demux_003_src22_valid),         //           .valid
		.src22_data          (cmd_xbar_demux_003_src22_data),          //           .data
		.src22_channel       (cmd_xbar_demux_003_src22_channel),       //           .channel
		.src22_startofpacket (cmd_xbar_demux_003_src22_startofpacket), //           .startofpacket
		.src22_endofpacket   (cmd_xbar_demux_003_src22_endofpacket),   //           .endofpacket
		.src23_ready         (cmd_xbar_demux_003_src23_ready),         //      src23.ready
		.src23_valid         (cmd_xbar_demux_003_src23_valid),         //           .valid
		.src23_data          (cmd_xbar_demux_003_src23_data),          //           .data
		.src23_channel       (cmd_xbar_demux_003_src23_channel),       //           .channel
		.src23_startofpacket (cmd_xbar_demux_003_src23_startofpacket), //           .startofpacket
		.src23_endofpacket   (cmd_xbar_demux_003_src23_endofpacket)    //           .endofpacket
	);

	nios2_cmd_xbar_demux_004 cmd_xbar_demux_004 (
		.clk                (nios_clk_clk),                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_004_src_ready),             //      sink.ready
		.sink_channel       (addr_router_004_src_channel),           //          .channel
		.sink_data          (addr_router_004_src_data),              //          .data
		.sink_startofpacket (addr_router_004_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_004_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_004_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_mux_021 cmd_xbar_mux_021 (
		.clk                 (altpll_0_c0_clk),                        //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_021_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_021_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_021_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_021_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_021_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_021_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_003_src15_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_003_src15_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_003_src15_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_003_src15_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_003_src15_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_003_src15_endofpacket),   //          .endofpacket
		.sink1_ready         (crosser_001_out_ready),                  //     sink1.ready
		.sink1_valid         (crosser_001_out_valid),                  //          .valid
		.sink1_channel       (crosser_001_out_channel),                //          .channel
		.sink1_data          (crosser_001_out_data),                   //          .data
		.sink1_startofpacket (crosser_001_out_startofpacket),          //          .startofpacket
		.sink1_endofpacket   (crosser_001_out_endofpacket)             //          .endofpacket
	);

	nios2_cmd_xbar_mux_021 cmd_xbar_mux_022 (
		.clk                 (altpll_0_c0_clk),                        //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_022_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_022_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_022_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_022_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_022_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_022_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_003_src16_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_003_src16_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_003_src16_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_003_src16_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_003_src16_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_003_src16_endofpacket),   //          .endofpacket
		.sink1_ready         (crosser_002_out_ready),                  //     sink1.ready
		.sink1_valid         (crosser_002_out_valid),                  //          .valid
		.sink1_channel       (crosser_002_out_channel),                //          .channel
		.sink1_data          (crosser_002_out_data),                   //          .data
		.sink1_startofpacket (crosser_002_out_startofpacket),          //          .startofpacket
		.sink1_endofpacket   (crosser_002_out_endofpacket)             //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_007 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_008 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_009 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_010 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_011 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_012 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_013 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_014 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_015 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_016 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_017 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_018 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_019 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_020 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_demux_004 rsp_xbar_demux_021 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_021_src_ready),               //      sink.ready
		.sink_channel       (id_router_021_src_channel),             //          .channel
		.sink_data          (id_router_021_src_data),                //          .data
		.sink_startofpacket (id_router_021_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_021_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_021_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_021_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_021_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_021_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_021_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_021_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_021_src1_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_demux_004 rsp_xbar_demux_022 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_022_src_ready),               //      sink.ready
		.sink_channel       (id_router_022_src_channel),             //          .channel
		.sink_data          (id_router_022_src_data),                //          .data
		.sink_startofpacket (id_router_022_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_022_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_022_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_022_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_022_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_022_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_022_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_022_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_022_src1_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_023 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_023_src_ready),               //      sink.ready
		.sink_channel       (id_router_023_src_channel),             //          .channel
		.sink_data          (id_router_023_src_data),                //          .data
		.sink_startofpacket (id_router_023_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_023_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_023_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_023_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_023_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_024 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_024_src_ready),               //      sink.ready
		.sink_channel       (id_router_024_src_channel),             //          .channel
		.sink_data          (id_router_024_src_data),                //          .data
		.sink_startofpacket (id_router_024_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_024_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_024_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_024_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_024_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_025 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_025_src_ready),               //      sink.ready
		.sink_channel       (id_router_025_src_channel),             //          .channel
		.sink_data          (id_router_025_src_data),                //          .data
		.sink_startofpacket (id_router_025_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_025_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_025_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_025_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_025_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_026 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_026_src_ready),               //      sink.ready
		.sink_channel       (id_router_026_src_channel),             //          .channel
		.sink_data          (id_router_026_src_data),                //          .data
		.sink_startofpacket (id_router_026_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_026_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_026_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_026_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_026_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_027 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_027_src_ready),               //      sink.ready
		.sink_channel       (id_router_027_src_channel),             //          .channel
		.sink_data          (id_router_027_src_data),                //          .data
		.sink_startofpacket (id_router_027_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_027_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_027_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_027_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_027_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_028 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_028_src_ready),               //      sink.ready
		.sink_channel       (id_router_028_src_channel),             //          .channel
		.sink_data          (id_router_028_src_data),                //          .data
		.sink_startofpacket (id_router_028_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_028_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_028_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_028_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_028_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_006 rsp_xbar_demux_029 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_029_src_ready),               //      sink.ready
		.sink_channel       (id_router_029_src_channel),             //          .channel
		.sink_data          (id_router_029_src_data),                //          .data
		.sink_startofpacket (id_router_029_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_029_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_029_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_029_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_029_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_mux_003 rsp_xbar_mux_003 (
		.clk                  (altpll_0_c0_clk),                       //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_003_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_003_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_003_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready          (crosser_003_out_ready),                 //     sink0.ready
		.sink0_valid          (crosser_003_out_valid),                 //          .valid
		.sink0_channel        (crosser_003_out_channel),               //          .channel
		.sink0_data           (crosser_003_out_data),                  //          .data
		.sink0_startofpacket  (crosser_003_out_startofpacket),         //          .startofpacket
		.sink0_endofpacket    (crosser_003_out_endofpacket),           //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_007_src0_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_008_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_009_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_010_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_010_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_011_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_011_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_012_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_012_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_013_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_013_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_014_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_014_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_015_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_015_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_016_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_017_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_018_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_019_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_020_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_021_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_022_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_023_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_024_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_024_src0_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_025_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_025_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_026_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_026_src0_endofpacket),   //          .endofpacket
		.sink21_ready         (rsp_xbar_demux_027_src0_ready),         //    sink21.ready
		.sink21_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.sink21_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.sink21_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.sink21_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.sink21_endofpacket   (rsp_xbar_demux_027_src0_endofpacket),   //          .endofpacket
		.sink22_ready         (rsp_xbar_demux_028_src0_ready),         //    sink22.ready
		.sink22_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.sink22_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.sink22_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.sink22_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.sink22_endofpacket   (rsp_xbar_demux_028_src0_endofpacket),   //          .endofpacket
		.sink23_ready         (rsp_xbar_demux_029_src0_ready),         //    sink23.ready
		.sink23_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.sink23_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.sink23_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.sink23_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.sink23_endofpacket   (rsp_xbar_demux_029_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_mux_004 rsp_xbar_mux_004 (
		.clk                 (nios_clk_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),     // clk_reset.reset
		.src_ready           (rsp_xbar_mux_004_src_ready),         //       src.ready
		.src_valid           (rsp_xbar_mux_004_src_valid),         //          .valid
		.src_data            (rsp_xbar_mux_004_src_data),          //          .data
		.src_channel         (rsp_xbar_mux_004_src_channel),       //          .channel
		.src_startofpacket   (rsp_xbar_mux_004_src_startofpacket), //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_004_src_endofpacket),   //          .endofpacket
		.sink0_ready         (crosser_004_out_ready),              //     sink0.ready
		.sink0_valid         (crosser_004_out_valid),              //          .valid
		.sink0_channel       (crosser_004_out_channel),            //          .channel
		.sink0_data          (crosser_004_out_data),               //          .data
		.sink0_startofpacket (crosser_004_out_startofpacket),      //          .startofpacket
		.sink0_endofpacket   (crosser_004_out_endofpacket),        //          .endofpacket
		.sink1_ready         (crosser_005_out_ready),              //     sink1.ready
		.sink1_valid         (crosser_005_out_valid),              //          .valid
		.sink1_channel       (crosser_005_out_channel),            //          .channel
		.sink1_data          (crosser_005_out_data),               //          .data
		.sink1_startofpacket (crosser_005_out_startofpacket),      //          .startofpacket
		.sink1_endofpacket   (crosser_005_out_endofpacket)         //          .endofpacket
	);

	nios2_cmd_xbar_demux_005 cmd_xbar_demux_005 (
		.clk                (ddr2_sysclk_clk),                       //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_005_src_ready),             //      sink.ready
		.sink_channel       (addr_router_005_src_channel),           //          .channel
		.sink_data          (addr_router_005_src_data),              //          .data
		.sink_startofpacket (addr_router_005_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_005_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_005_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_demux_005 rsp_xbar_demux_030 (
		.clk                (ddr2_sysclk_clk),                       //       clk.clk
		.reset              (~ddr2_reset_request_n_reset),           // clk_reset.reset
		.sink_ready         (id_router_030_src_ready),               //      sink.ready
		.sink_channel       (id_router_030_src_channel),             //          .channel
		.sink_data          (id_router_030_src_data),                //          .data
		.sink_startofpacket (id_router_030_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_030_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_030_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_030_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_030_src0_endofpacket)    //          .endofpacket
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (85),
		.BITS_PER_SYMBOL     (85),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (24),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (altpll_0_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_004_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_003_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_003_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_003_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_003_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_003_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_003_src0_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (85),
		.BITS_PER_SYMBOL     (85),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (24),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (nios_clk_clk),                          //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (altpll_0_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (85),
		.BITS_PER_SYMBOL     (85),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (24),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (nios_clk_clk),                          //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (altpll_0_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src1_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src1_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src1_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src1_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src1_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src1_data),          //              .data
		.out_ready         (crosser_002_out_ready),                 //           out.ready
		.out_valid         (crosser_002_out_valid),                 //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_002_out_channel),               //              .channel
		.out_data          (crosser_002_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (85),
		.BITS_PER_SYMBOL     (85),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (24),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_004_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_006_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_006_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_006_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_006_src0_data),          //              .data
		.out_ready         (crosser_003_out_ready),                 //           out.ready
		.out_valid         (crosser_003_out_valid),                 //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_003_out_channel),               //              .channel
		.out_data          (crosser_003_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (85),
		.BITS_PER_SYMBOL     (85),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (24),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_004 (
		.in_clk            (altpll_0_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (nios_clk_clk),                          //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_021_src1_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_021_src1_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_021_src1_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_021_src1_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_021_src1_channel),       //              .channel
		.in_data           (rsp_xbar_demux_021_src1_data),          //              .data
		.out_ready         (crosser_004_out_ready),                 //           out.ready
		.out_valid         (crosser_004_out_valid),                 //              .valid
		.out_startofpacket (crosser_004_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_004_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_004_out_channel),               //              .channel
		.out_data          (crosser_004_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (85),
		.BITS_PER_SYMBOL     (85),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (24),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_005 (
		.in_clk            (altpll_0_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (nios_clk_clk),                          //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_022_src1_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_022_src1_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_022_src1_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_022_src1_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_022_src1_channel),       //              .channel
		.in_data           (rsp_xbar_demux_022_src1_data),          //              .data
		.out_ready         (crosser_005_out_ready),                 //           out.ready
		.out_valid         (crosser_005_out_valid),                 //              .valid
		.out_startofpacket (crosser_005_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_005_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_005_out_channel),               //              .channel
		.out_data          (crosser_005_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	nios2_irq_mapper irq_mapper (
		.clk            (nios_clk_clk),                   //        clk.clk
		.reset          (rst_controller_reset_out_reset), //  clk_reset.reset
		.receiver0_irq  (irq_mapper_receiver0_irq),       //  receiver0.irq
		.receiver1_irq  (irq_mapper_receiver1_irq),       //  receiver1.irq
		.receiver2_irq  (irq_mapper_receiver2_irq),       //  receiver2.irq
		.receiver3_irq  (irq_mapper_receiver3_irq),       //  receiver3.irq
		.receiver4_irq  (irq_mapper_receiver4_irq),       //  receiver4.irq
		.receiver5_irq  (irq_mapper_receiver5_irq),       //  receiver5.irq
		.receiver6_irq  (irq_mapper_receiver6_irq),       //  receiver6.irq
		.receiver7_irq  (irq_mapper_receiver7_irq),       //  receiver7.irq
		.receiver8_irq  (irq_mapper_receiver8_irq),       //  receiver8.irq
		.receiver9_irq  (irq_mapper_receiver9_irq),       //  receiver9.irq
		.receiver10_irq (irq_mapper_receiver10_irq),      // receiver10.irq
		.receiver11_irq (irq_mapper_receiver11_irq),      // receiver11.irq
		.sender_irq     (nios2_d_irq_irq)                 //     sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_0_c0_clk),                    //       receiver_clk.clk
		.sender_clk     (nios_clk_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (altpll_0_c0_clk),                    //       receiver_clk.clk
		.sender_clk     (nios_clk_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (altpll_0_c0_clk),                    //       receiver_clk.clk
		.sender_clk     (nios_clk_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (altpll_0_c0_clk),                    //       receiver_clk.clk
		.sender_clk     (nios_clk_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (altpll_0_c0_clk),                    //       receiver_clk.clk
		.sender_clk     (nios_clk_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_005 (
		.receiver_clk   (altpll_0_c0_clk),                    //       receiver_clk.clk
		.sender_clk     (nios_clk_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_005_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver7_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_006 (
		.receiver_clk   (altpll_0_c0_clk),                    //       receiver_clk.clk
		.sender_clk     (nios_clk_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_006_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver8_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_007 (
		.receiver_clk   (altpll_0_c0_clk),                    //       receiver_clk.clk
		.sender_clk     (nios_clk_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_007_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver9_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_008 (
		.receiver_clk   (altpll_0_c0_clk),                    //       receiver_clk.clk
		.sender_clk     (nios_clk_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_008_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver10_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_009 (
		.receiver_clk   (altpll_0_c0_clk),                    //       receiver_clk.clk
		.sender_clk     (nios_clk_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_009_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver11_irq)           //             sender.irq
	);

endmodule
